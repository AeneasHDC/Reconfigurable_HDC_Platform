----
 -- @file level_hvec_gen_hdl.hpp
 -- @brief This script generates HDL code for generating high-dimensional LEVEL vectors.
 -- It is a novel method; for more information, please refer to our paper.
 --
 -- @author Saeid Jamili and Marco Angioli
 -- @note Author names are listed in alphabetical order.
 -- @email <saeid.jamili@uniroma1.it>
 -- @email <marco.angioli@uniroma1.it>
 --
 -- @contributors
 --
 -- @date Created: 24th July 2023
 -- @date Last Updated: 23th August 2023
 --
 -- @version 1.0.0
 --
 -- @institute Sapienza University of Rome
 -- @cite https://doi.org/10.xxxx/yyyyy
 --
 -- @section DEPENDENCIES
 -- - Dependency1: Description or version details.
 -- - Dependency2: Description or version details.
 --
 -- @section LICENSE
 -- This file is part of the Aeneas HyperCompute Platform.
 --
 -- Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 --
 -- @section CHANGELOG
 -- @version 1.0.0-dev - 23th August 2023
 -- - Initial release
 --
 -- @todo
 -- - Complete level vector generator function
 -- - Add training
 --
 -- @see
 -- -
 -- -
 -- -
 --
 --

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity level_vec_gen is
    Port ( level_vec_out : out  STD_LOGIC_VECTOR (63 downto 0);
           frame_index : in  STD_LOGIC_VECTOR (2 downto 0);
           frame_id : in  STD_LOGIC_VECTOR (4 downto 0));
end level_vec_gen;

architecture Behavioral of level_vec_gen is
begin
    process (frame_index, frame_id)
    begin
        -- Update this function to match your requirements
        case frame_index is
            when "000" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1111100011110101011011110101100111100000010100101000101000110000";
                    when "00001" => level_vec_out <= "1111100011110101011011110101100111100000010100101000101000110000";
                    when "00010" => level_vec_out <= "1111101011110101011011110101100111100000010100101000101000110000";
                    when "00011" => level_vec_out <= "1111101011110101011011110101100111100000010100101000101000110000";
                    when "00100" => level_vec_out <= "1111101011110101011011110101100111100000010100101000101000110000";
                    when "00101" => level_vec_out <= "1111101011111101011011110101100111100010010100101000101000110000";
                    when "00110" => level_vec_out <= "1111101011111101011011110101100111100010010101101000101000110000";
                    when "00111" => level_vec_out <= "1111101011111101011011110101100111100010011101101000101000110000";
                    when "01000" => level_vec_out <= "1111101011111101011011110101100111100010011101101000101000110000";
                    when "01001" => level_vec_out <= "1111101011111101011011110101110111100010011101101000101000110000";
                    when "01010" => level_vec_out <= "1111101011111101011011110101111111100011111101101000101000110000";
                    when "01011" => level_vec_out <= "1111101011111101011011110101111111100011111101101000111000110001";
                    when "01100" => level_vec_out <= "1111101011111101011111110101111111100011111101101000111000110001";
                    when "01101" => level_vec_out <= "1111101011111101011111110101111111100011111101101000111000110001";
                    when "01110" => level_vec_out <= "1111101011111101011111110101111111100011111101101000111000111011";
                    when "01111" => level_vec_out <= "1111101011111101011111110101111111100011111101101000111100111011";
                    when "10000" => level_vec_out <= "1111101011111101011111110101111111100011111101101000111100111011";
                    when "10001" => level_vec_out <= "1111101011111111011111110101111111100011111101101000111100111011";
                    when "10010" => level_vec_out <= "1111101011111111011111110101111111100011111101101000111100111011";
                    when "10011" => level_vec_out <= "1111101011111111011111110101111111100011111101101001111100111011";
                    when "10100" => level_vec_out <= "1111101011111111011111110101111111100011111101101001111101111011";
                    when "10101" => level_vec_out <= "1111101011111111011111110101111111111011111101101101111101111011";
                    when "10110" => level_vec_out <= "1111101011111111011111110101111111111011111101101101111101111111";
                    when "10111" => level_vec_out <= "1111101011111111011111110101111111111011111101101101111101111111";
                    when "11000" => level_vec_out <= "1111101011111111011111111101111111111111111101101101111101111111";
                    when "11001" => level_vec_out <= "1111101011111111011111111101111111111111111101101101111101111111";
                    when "11010" => level_vec_out <= "1111101011111111011111111101111111111111111101111101111101111111";
                    when "11011" => level_vec_out <= "1111101011111111111111111101111111111111111101111101111101111111";
                    when "11100" => level_vec_out <= "1111101011111111111111111101111111111111111101111101111111111111";
                    when "11101" => level_vec_out <= "1111101011111111111111111111111111111111111101111101111111111111";
                    when "11110" => level_vec_out <= "1111111011111111111111111111111111111111111101111101111111111111";
                    when "11111" => level_vec_out <= "1111111011111111111111111111111111111111111101111111111111111111";
                when others => null;
                end case;
            when "001" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1010100001101100010010010010110000011001000010000000001111011111";
                    when "00001" => level_vec_out <= "1010100001101100010010010010110000011001000010100000001111011111";
                    when "00010" => level_vec_out <= "1010100001101100010011010010110000011001000010100000001111011111";
                    when "00011" => level_vec_out <= "1010100001101100010111010010110000011001000010100000001111011111";
                    when "00100" => level_vec_out <= "1110100001101110010111010010110000011001001010100000001111011111";
                    when "00101" => level_vec_out <= "1110100101101111010111010010110100011001001010100000001111011111";
                    when "00110" => level_vec_out <= "1110100101101111010111010010110100011001001010100000101111011111";
                    when "00111" => level_vec_out <= "1110100101101111010111010010110100011001001010100000101111011111";
                    when "01000" => level_vec_out <= "1110100101101111011111010010110100011001001010100000101111011111";
                    when "01001" => level_vec_out <= "1110100101101111011111010010111100011001001010100000101111011111";
                    when "01010" => level_vec_out <= "1110100101101111011111010010111100011001001010100010101111011111";
                    when "01011" => level_vec_out <= "1110100101101111011111010010111100011001001010100011101111011111";
                    when "01100" => level_vec_out <= "1110100111101111011111010011111100011001001010100011101111011111";
                    when "01101" => level_vec_out <= "1110100111101111011111010011111100011001011010110011101111011111";
                    when "01110" => level_vec_out <= "1110100111101111011111010011111100011001011010110011101111011111";
                    when "01111" => level_vec_out <= "1110100111101111011111010011111100011001011010110011101111011111";
                    when "10000" => level_vec_out <= "1110100111101111011111010011111100011011011010110111101111011111";
                    when "10001" => level_vec_out <= "1110100111101111011111010011111100011011011010110111101111011111";
                    when "10010" => level_vec_out <= "1110101111101111011111010011111100011011011011110111111111011111";
                    when "10011" => level_vec_out <= "1110101111101111011111010011111100011011011011110111111111011111";
                    when "10100" => level_vec_out <= "1110101111101111111111010111111100011011011011110111111111011111";
                    when "10101" => level_vec_out <= "1110101111111111111111010111111100011011011111111111111111011111";
                    when "10110" => level_vec_out <= "1110101111111111111111011111111100011011011111111111111111011111";
                    when "10111" => level_vec_out <= "1111101111111111111111011111111100011011011111111111111111011111";
                    when "11000" => level_vec_out <= "1111101111111111111111011111111100111011011111111111111111011111";
                    when "11001" => level_vec_out <= "1111101111111111111111011111111100111011011111111111111111111111";
                    when "11010" => level_vec_out <= "1111111111111111111111011111111100111011011111111111111111111111";
                    when "11011" => level_vec_out <= "1111111111111111111111011111111100111111011111111111111111111111";
                    when "11100" => level_vec_out <= "1111111111111111111111011111111101111111011111111111111111111111";
                    when "11101" => level_vec_out <= "1111111111111111111111111111111111111111011111111111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111011111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "010" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0000010100010110010111010110110110001110110100010110110110010100";
                    when "00001" => level_vec_out <= "0000010100010110010111010110110110001110110110010110110110010100";
                    when "00010" => level_vec_out <= "0000010100010110010111010110110110001110110110010110110110010100";
                    when "00011" => level_vec_out <= "0000010100010110011111010110110110001110110110010110110110010100";
                    when "00100" => level_vec_out <= "0100010100010110011111010110110110001110110110010110110110010110";
                    when "00101" => level_vec_out <= "0100010100010110011111010110110110001110110110010110110110010110";
                    when "00110" => level_vec_out <= "0100010100010110011111010110110110001110110110011110110110010110";
                    when "00111" => level_vec_out <= "0100010100010111011111010110110110001110110110011110110110010110";
                    when "01000" => level_vec_out <= "0100010100010111011111011110110111001110110110011110110110010110";
                    when "01001" => level_vec_out <= "0100010100010111011111011110110111001110110111011110110110010110";
                    when "01010" => level_vec_out <= "0100010100010111011111011110110111001110110111011110110110010110";
                    when "01011" => level_vec_out <= "0100010100010111011111011110110111001110110111011110110110010111";
                    when "01100" => level_vec_out <= "0100010100010111011111011110110111001110110111011110110110010111";
                    when "01101" => level_vec_out <= "0100010100010111111111011110110111101110110111011110110110010111";
                    when "01110" => level_vec_out <= "0100010100010111111111011110110111101110110111011110110111010111";
                    when "01111" => level_vec_out <= "0110010100010111111111011110110111101111110111011110110111010111";
                    when "10000" => level_vec_out <= "0110010100010111111111111110110111101111110111011110110111010111";
                    when "10001" => level_vec_out <= "0110010100010111111111111110110111111111110111011110110111010111";
                    when "10010" => level_vec_out <= "0110010100010111111111111111110111111111110111011110110111010111";
                    when "10011" => level_vec_out <= "0110010100010111111111111111110111111111110111011110110111110111";
                    when "10100" => level_vec_out <= "0110010100010111111111111111110111111111110111011110110111110111";
                    when "10101" => level_vec_out <= "0110010100010111111111111111110111111111110111011110110111110111";
                    when "10110" => level_vec_out <= "0110010100010111111111111111110111111111110111011110110111110111";
                    when "10111" => level_vec_out <= "1110010100010111111111111111110111111111110111011110110111110111";
                    when "11000" => level_vec_out <= "1110010100010111111111111111110111111111110111111110110111110111";
                    when "11001" => level_vec_out <= "1110010100010111111111111111110111111111111111111111110111110111";
                    when "11010" => level_vec_out <= "1110010100010111111111111111110111111111111111111111110111110111";
                    when "11011" => level_vec_out <= "1110111100010111111111111111110111111111111111111111110111110111";
                    when "11100" => level_vec_out <= "1111111100011111111111111111110111111111111111111111110111110111";
                    when "11101" => level_vec_out <= "1111111100011111111111111111110111111111111111111111110111110111";
                    when "11110" => level_vec_out <= "1111111110111111111111111111110111111111111111111111110111110111";
                    when "11111" => level_vec_out <= "1111111110111111111111111111111111111111111111111111110111111111";
                when others => null;
                end case;
            when "011" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1011111001111111101000100111010001101100001001011000010000111110";
                    when "00001" => level_vec_out <= "1011111001111111111000100111010001101100101001011000010000111110";
                    when "00010" => level_vec_out <= "1011111001111111111000100111010001101100101001011000010000111110";
                    when "00011" => level_vec_out <= "1011111001111111111000100111010001101100101011011000010000111110";
                    when "00100" => level_vec_out <= "1011111001111111111000100111010001101100101011011000010000111110";
                    when "00101" => level_vec_out <= "1011111001111111111001100111010001101100101011011000010011111110";
                    when "00110" => level_vec_out <= "1011111001111111111001100111110001101100101011011000010011111110";
                    when "00111" => level_vec_out <= "1011111101111111111011100111110101101100101011011000010011111110";
                    when "01000" => level_vec_out <= "1011111101111111111011100111110101101110101011011101010011111110";
                    when "01001" => level_vec_out <= "1111111101111111111011100111110101101110101011011101010011111110";
                    when "01010" => level_vec_out <= "1111111111111111111011100111110101101110101011011101010111111110";
                    when "01011" => level_vec_out <= "1111111111111111111011100111110101101110101011011101010111111110";
                    when "01100" => level_vec_out <= "1111111111111111111011100111110101101110101011011101110111111110";
                    when "01101" => level_vec_out <= "1111111111111111111011100111110101101110101011011101110111111111";
                    when "01110" => level_vec_out <= "1111111111111111111011100111110101101110101111011101110111111111";
                    when "01111" => level_vec_out <= "1111111111111111111011100111110101101110101111011101110111111111";
                    when "10000" => level_vec_out <= "1111111111111111111011100111110101101110101111011101110111111111";
                    when "10001" => level_vec_out <= "1111111111111111111011100111110101101110101111011101110111111111";
                    when "10010" => level_vec_out <= "1111111111111111111011100111110101101110101111011101110111111111";
                    when "10011" => level_vec_out <= "1111111111111111111011100111110111101110101111011101110111111111";
                    when "10100" => level_vec_out <= "1111111111111111111011100111110111101110101111011101111111111111";
                    when "10101" => level_vec_out <= "1111111111111111111011100111110111101110101111011101111111111111";
                    when "10110" => level_vec_out <= "1111111111111111111011100111110111101110101111011101111111111111";
                    when "10111" => level_vec_out <= "1111111111111111111011110111110111101110101111011101111111111111";
                    when "11000" => level_vec_out <= "1111111111111111111011111111110111101110101111011101111111111111";
                    when "11001" => level_vec_out <= "1111111111111111111011111111110111101110111111011101111111111111";
                    when "11010" => level_vec_out <= "1111111111111111111011111111111111101111111111011111111111111111";
                    when "11011" => level_vec_out <= "1111111111111111111011111111111111101111111111011111111111111111";
                    when "11100" => level_vec_out <= "1111111111111111111011111111111111101111111111111111111111111111";
                    when "11101" => level_vec_out <= "1111111111111111111011111111111111101111111111111111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111011111111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111011111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "100" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1001110001111110111000000100000111101110110001010111010010010100";
                    when "00001" => level_vec_out <= "1001110001111110111000000110000111101110110001110111010010010100";
                    when "00010" => level_vec_out <= "1001110001111110111000000110000111101110110001110111010010010100";
                    when "00011" => level_vec_out <= "1011110001111110111000000110000111101110110001110111010010010100";
                    when "00100" => level_vec_out <= "1011110001111110111000000110000111101110110001110111010010010100";
                    when "00101" => level_vec_out <= "1011110001111110111000000110000111101110110001110111010010010100";
                    when "00110" => level_vec_out <= "1111110001111110111000000111000111101110110001110111010010010100";
                    when "00111" => level_vec_out <= "1111110001111110111000000111000111101110111001110111010010010100";
                    when "01000" => level_vec_out <= "1111110001111110111000000111000111101110111001110111010010010100";
                    when "01001" => level_vec_out <= "1111110001111110111000000111000111101110111001110111010010010100";
                    when "01010" => level_vec_out <= "1111110001111110111000000111000111101110111001110111010010010100";
                    when "01011" => level_vec_out <= "1111110001111110111000000111000111101110111001110111010010010100";
                    when "01100" => level_vec_out <= "1111110001111110111000000111000111101110111001110111010010010100";
                    when "01101" => level_vec_out <= "1111110001111110111000000111000111101110111001110111010010010100";
                    when "01110" => level_vec_out <= "1111110001111110111001000111000111101110111001111111010010010100";
                    when "01111" => level_vec_out <= "1111110001111110111001101111000111101110111001111111010011110100";
                    when "10000" => level_vec_out <= "1111110001111110111001101111010111101110111001111111010011110100";
                    when "10001" => level_vec_out <= "1111110001111110111001101111010111101110111011111111011011110100";
                    when "10010" => level_vec_out <= "1111110001111110111011101111010111101110111111111111011111110100";
                    when "10011" => level_vec_out <= "1111110001111111111011101111010111101111111111111111011111110100";
                    when "10100" => level_vec_out <= "1111110001111111111111101111011111101111111111111111011111110100";
                    when "10101" => level_vec_out <= "1111110001111111111111101111011111101111111111111111011111110100";
                    when "10110" => level_vec_out <= "1111111011111111111111111111011111101111111111111111011111110100";
                    when "10111" => level_vec_out <= "1111111011111111111111111111011111101111111111111111011111111100";
                    when "11000" => level_vec_out <= "1111111011111111111111111111111111101111111111111111011111111101";
                    when "11001" => level_vec_out <= "1111111011111111111111111111111111101111111111111111011111111101";
                    when "11010" => level_vec_out <= "1111111011111111111111111111111111101111111111111111011111111111";
                    when "11011" => level_vec_out <= "1111111011111111111111111111111111111111111111111111011111111111";
                    when "11100" => level_vec_out <= "1111111011111111111111111111111111111111111111111111111111111111";
                    when "11101" => level_vec_out <= "1111111011111111111111111111111111111111111111111111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "101" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0101011101100111110101010111110110100111100011111010101010101111";
                    when "00001" => level_vec_out <= "0101011101100111110101010111110110100111100011111010101010101111";
                    when "00010" => level_vec_out <= "0101011101100111110111010111110110100111100011111010101010101111";
                    when "00011" => level_vec_out <= "0101011101100111110111010111110110100111100011111011101011101111";
                    when "00100" => level_vec_out <= "1101011101100111110111010111110111100111100011111011101011101111";
                    when "00101" => level_vec_out <= "1101011101100111110111010111110111100111100011111011101011101111";
                    when "00110" => level_vec_out <= "1101011101100111110111010111110111100111100011111011101011101111";
                    when "00111" => level_vec_out <= "1101011101100111110111010111110111100111100011111011101011101111";
                    when "01000" => level_vec_out <= "1101011101100111110111010111110111100111100011111011101011101111";
                    when "01001" => level_vec_out <= "1101011101100111110111010111110111100111100011111011101011101111";
                    when "01010" => level_vec_out <= "1101011101100111110111010111110111100111110011111011101011101111";
                    when "01011" => level_vec_out <= "1101011101100111111111010111110111100111110011111011111011101111";
                    when "01100" => level_vec_out <= "1101011101100111111111110111110111101111110011111111111011101111";
                    when "01101" => level_vec_out <= "1101011101100111111111110111110111101111110011111111111011101111";
                    when "01110" => level_vec_out <= "1101011101100111111111110111110111101111110011111111111011101111";
                    when "01111" => level_vec_out <= "1101011101100111111111110111110111101111110011111111111011101111";
                    when "10000" => level_vec_out <= "1101111101101111111111110111110111101111110011111111111011101111";
                    when "10001" => level_vec_out <= "1101111101101111111111110111110111101111110011111111111011101111";
                    when "10010" => level_vec_out <= "1101111101101111111111110111110111101111110011111111111011101111";
                    when "10011" => level_vec_out <= "1101111101101111111111110111110111101111110111111111111011101111";
                    when "10100" => level_vec_out <= "1101111101101111111111110111110111101111110111111111111011101111";
                    when "10101" => level_vec_out <= "1101111101101111111111110111110111101111110111111111111011101111";
                    when "10110" => level_vec_out <= "1101111101101111111111110111110111101111110111111111111011111111";
                    when "10111" => level_vec_out <= "1101111101101111111111110111110111101111110111111111111011111111";
                    when "11000" => level_vec_out <= "1101111101101111111111111111110111101111110111111111111011111111";
                    when "11001" => level_vec_out <= "1101111101101111111111111111110111101111110111111111111011111111";
                    when "11010" => level_vec_out <= "1101111101111111111111111111110111101111110111111111111011111111";
                    when "11011" => level_vec_out <= "1101111101111111111111111111110111111111110111111111111011111111";
                    when "11100" => level_vec_out <= "1101111101111111111111111111110111111111110111111111111011111111";
                    when "11101" => level_vec_out <= "1101111111111111111111111111110111111111111111111111111011111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111110111111111111111111111111011111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "110" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0110000011000110001100101111110000100110001101001010100100000001";
                    when "00001" => level_vec_out <= "0110000011000110001100101111110000100110101101001010100100000001";
                    when "00010" => level_vec_out <= "0111000011001110001100101111110000100110101101001010100100000001";
                    when "00011" => level_vec_out <= "0111000011001110001100101111110001100110101101001010100100000001";
                    when "00100" => level_vec_out <= "0111000011001110001100101111110001100110101101001010100100000001";
                    when "00101" => level_vec_out <= "0111000011001110001100101111110001100110101101001010100100000001";
                    when "00110" => level_vec_out <= "0111000111001110001100101111110001100110101101001010100100000001";
                    when "00111" => level_vec_out <= "0111000111001110001100101111110001100110101101001010110101000001";
                    when "01000" => level_vec_out <= "0111000111001110001100101111110001100110101101001010110101000001";
                    when "01001" => level_vec_out <= "0111000111001110001100101111110011100110101101001010110101000001";
                    when "01010" => level_vec_out <= "0111000111001110001100101111110011100110101101001110110101000001";
                    when "01011" => level_vec_out <= "0111011111001110001100101111110011100110101101001110110101000001";
                    when "01100" => level_vec_out <= "0111011111001110001100101111110111100110101101001110110101000001";
                    when "01101" => level_vec_out <= "1111011111001110001100101111111111100110101101001110110101000001";
                    when "01110" => level_vec_out <= "1111011111001110001100101111111111100110101101001110110101000011";
                    when "01111" => level_vec_out <= "1111011111001110001100101111111111100110101101001110110101000011";
                    when "10000" => level_vec_out <= "1111011111001110001101101111111111100110101101001110110101000011";
                    when "10001" => level_vec_out <= "1111011111001110001101101111111111100110101101001110111101000111";
                    when "10010" => level_vec_out <= "1111011111001110001101101111111111100110101101001110111101000111";
                    when "10011" => level_vec_out <= "1111011111011110001101101111111111100110101101001110111101000111";
                    when "10100" => level_vec_out <= "1111011111111110001101101111111111100110111101001110111101000111";
                    when "10101" => level_vec_out <= "1111011111111110001101101111111111101110111101001110111101000111";
                    when "10110" => level_vec_out <= "1111011111111110001101101111111111101110111101001110111101001111";
                    when "10111" => level_vec_out <= "1111011111111110111101101111111111101110111101001111111101001111";
                    when "11000" => level_vec_out <= "1111011111111110111101101111111111101110111101001111111101001111";
                    when "11001" => level_vec_out <= "1111011111111111111101101111111111111110111111001111111101001111";
                    when "11010" => level_vec_out <= "1111111111111111111101101111111111111110111111001111111101001111";
                    when "11011" => level_vec_out <= "1111111111111111111101111111111111111110111111011111111101001111";
                    when "11100" => level_vec_out <= "1111111111111111111101111111111111111110111111011111111101101111";
                    when "11101" => level_vec_out <= "1111111111111111111101111111111111111110111111111111111101111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111110111111111111111101111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111110111111111111111101111111";
                when others => null;
                end case;
            when "111" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1110010101010110011111010001010100111000101001111110100011001010";
                    when "00001" => level_vec_out <= "1110010101010110011111010001010100111000101001111110110011001010";
                    when "00010" => level_vec_out <= "1110010101010110011111010011010100111010111001111110110011001010";
                    when "00011" => level_vec_out <= "1110010101010110011111010011010100111010111011111110110011001010";
                    when "00100" => level_vec_out <= "1110010101010110011111010011010100111110111011111110110011001010";
                    when "00101" => level_vec_out <= "1110010101010110011111010011010100111110111011111110110011001010";
                    when "00110" => level_vec_out <= "1110010101010110011111010011010100111110111011111110111011001010";
                    when "00111" => level_vec_out <= "1110010101010110011111010011010100111110111011111110111011001010";
                    when "01000" => level_vec_out <= "1110011101011110011111010011010100111110111011111110111011001010";
                    when "01001" => level_vec_out <= "1110011101011111011111010111010100111111111011111110111011001010";
                    when "01010" => level_vec_out <= "1110011101011111011111010111010100111111111011111110111011001010";
                    when "01011" => level_vec_out <= "1110011101011111011111010111010100111111111011111110111011001010";
                    when "01100" => level_vec_out <= "1110011101011111011111010111010100111111111011111110111011001010";
                    when "01101" => level_vec_out <= "1110011101011111011111010111010100111111111011111110111011011010";
                    when "01110" => level_vec_out <= "1110011101011111011111010111010100111111111011111110111111011010";
                    when "01111" => level_vec_out <= "1110011101011111011111010111010100111111111011111110111111111010";
                    when "10000" => level_vec_out <= "1110111101011111011111010111010100111111111011111110111111111010";
                    when "10001" => level_vec_out <= "1110111101011111011111010111011110111111111011111110111111111010";
                    when "10010" => level_vec_out <= "1110111101011111111111010111011110111111111011111110111111111010";
                    when "10011" => level_vec_out <= "1110111101011111111111010111011110111111111011111111111111111010";
                    when "10100" => level_vec_out <= "1110111101011111111111010111011110111111111011111111111111111010";
                    when "10101" => level_vec_out <= "1111111101011111111111010111011110111111111011111111111111111010";
                    when "10110" => level_vec_out <= "1111111101011111111111010111111110111111111011111111111111111010";
                    when "10111" => level_vec_out <= "1111111101011111111111010111111111111111111011111111111111111010";
                    when "11000" => level_vec_out <= "1111111101011111111111010111111111111111111011111111111111111010";
                    when "11001" => level_vec_out <= "1111111101011111111111010111111111111111111011111111111111111011";
                    when "11010" => level_vec_out <= "1111111101011111111111010111111111111111111011111111111111111011";
                    when "11011" => level_vec_out <= "1111111101011111111111010111111111111111111011111111111111111011";
                    when "11100" => level_vec_out <= "1111111101011111111111010111111111111111111111111111111111111011";
                    when "11101" => level_vec_out <= "1111111101011111111111110111111111111111111111111111111111111011";
                    when "11110" => level_vec_out <= "1111111111011111111111110111111111111111111111111111111111111011";
                    when "11111" => level_vec_out <= "1111111111011111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when others => null;
        end case;
    end process;
end Behavioral;