----
 -- @file level_hvec_gen_hdl.hpp
 -- @brief This script generates HDL code for generating high-dimensional LEVEL vectors.
 -- It is a novel method; for more information, please refer to our paper.
 --
 -- @author Saeid Jamili and Marco Angioli
 -- @note Author names are listed in alphabetical order.
 -- @email <saeid.jamili@uniroma1.it>
 -- @email <marco.angioli@uniroma1.it>
 --
 -- @contributors
 --
 -- @date Created: 24th July 2023
 -- @date Last Updated: 23th August 2023
 --
 -- @version 1.0.0
 --
 -- @institute Sapienza University of Rome
 -- @cite https://doi.org/10.xxxx/yyyyy
 --
 -- @section DEPENDENCIES
 -- - Dependency1: Description or version details.
 -- - Dependency2: Description or version details.
 --
 -- @section LICENSE
 -- This file is part of the Aeneas HyperCompute Platform.
 --
 -- Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 --
 -- @section CHANGELOG
 -- @version 1.0.0-dev - 23th August 2023
 -- - Initial release
 --
 -- @todo
 -- - Complete level vector generator function
 -- - Add training
 --
 -- @see
 -- -
 -- -
 -- -
 --
 --

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity level_vec_gen is
    Port ( level_vec_out : out  STD_LOGIC_VECTOR (63 downto 0);
           frame_index : in  STD_LOGIC_VECTOR (2 downto 0);
           frame_id : in  STD_LOGIC_VECTOR (4 downto 0));
end level_vec_gen;

architecture Behavioral of level_vec_gen is
begin
    process (frame_index, frame_id)
    begin
        -- Update this function to match your requirements
        case frame_index is
            when "000" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1110100110111100001011010111110100011111010000010010010001111111";
                    when "00001" => level_vec_out <= "1110100110111110011011110111110100011111010000010010010001111111";
                    when "00010" => level_vec_out <= "1110100110111110011011110111110100011111010000010110010001111111";
                    when "00011" => level_vec_out <= "1110100110111110011111110111110100011111010000010111010001111111";
                    when "00100" => level_vec_out <= "1110100110111110011111110111110100011111010000010111010001111111";
                    when "00101" => level_vec_out <= "1110100110111111011111110111111100011111010000010111010001111111";
                    when "00110" => level_vec_out <= "1110100110111111011111110111111100011111010000010111010011111111";
                    when "00111" => level_vec_out <= "1110100110111111011111110111111100111111010000010111010011111111";
                    when "01000" => level_vec_out <= "1110100110111111011111110111111100111111010000010111010011111111";
                    when "01001" => level_vec_out <= "1110100110111111011111110111111100111111010000010111010011111111";
                    when "01010" => level_vec_out <= "1110100110111111011111110111111100111111010000010111010011111111";
                    when "01011" => level_vec_out <= "1110100110111111011111110111111100111111010000010111010011111111";
                    when "01100" => level_vec_out <= "1110100110111111111111110111111100111111010000010111010011111111";
                    when "01101" => level_vec_out <= "1110100110111111111111110111111100111111010000010111010011111111";
                    when "01110" => level_vec_out <= "1110100110111111111111110111111100111111010000010111010111111111";
                    when "01111" => level_vec_out <= "1110100110111111111111110111111100111111010000010111010111111111";
                    when "10000" => level_vec_out <= "1110100110111111111111110111111101111111010000010111010111111111";
                    when "10001" => level_vec_out <= "1110100110111111111111110111111101111111010000010111010111111111";
                    when "10010" => level_vec_out <= "1110100110111111111111110111111101111111010000010111010111111111";
                    when "10011" => level_vec_out <= "1110100110111111111111110111111101111111110010010111010111111111";
                    when "10100" => level_vec_out <= "1110100110111111111111110111111101111111110010010111010111111111";
                    when "10101" => level_vec_out <= "1110100110111111111111110111111101111111110110010111010111111111";
                    when "10110" => level_vec_out <= "1110100110111111111111110111111101111111110110010111010111111111";
                    when "10111" => level_vec_out <= "1110100110111111111111110111111101111111110110010111010111111111";
                    when "11000" => level_vec_out <= "1110100110111111111111110111111101111111110110010111110111111111";
                    when "11001" => level_vec_out <= "1110101111111111111111110111111101111111110111010111110111111111";
                    when "11010" => level_vec_out <= "1110101111111111111111110111111101111111110111010111110111111111";
                    when "11011" => level_vec_out <= "1110101111111111111111110111111101111111110111010111110111111111";
                    when "11100" => level_vec_out <= "1110101111111111111111110111111111111111110111010111110111111111";
                    when "11101" => level_vec_out <= "1110101111111111111111111111111111111111110111010111110111111111";
                    when "11110" => level_vec_out <= "1111101111111111111111111111111111111111111111011111110111111111";
                    when "11111" => level_vec_out <= "1111101111111111111111111111111111111111111111111111110111111111";
                when others => null;
                end case;
            when "001" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1001000000101100111000110100010000111010010000001001111001100101";
                    when "00001" => level_vec_out <= "1001000000101100111000110100010000111010010000001001111001100101";
                    when "00010" => level_vec_out <= "1001000000101100111000110100010000111010010000001001111001100101";
                    when "00011" => level_vec_out <= "1001100000101100111000110100010000111010010001001001111001100101";
                    when "00100" => level_vec_out <= "1001100000101100111000110100011011111010010001001001111001101101";
                    when "00101" => level_vec_out <= "1001100000101101111000110100011011111010010001001001111001101101";
                    when "00110" => level_vec_out <= "1001100000101101111010110100011011111010010001001001111001101101";
                    when "00111" => level_vec_out <= "1001101000101101111010110100011011111010010001001001111011101101";
                    when "01000" => level_vec_out <= "1001101000101101111010110101011011111010010001001001111011101101";
                    when "01001" => level_vec_out <= "1001101011101101111010110101011011111010010001001001111011101101";
                    when "01010" => level_vec_out <= "1001101011101101111010110101011011111010010001001001111011101101";
                    when "01011" => level_vec_out <= "1001101011111101111010110101011011111010010001001001111011101101";
                    when "01100" => level_vec_out <= "1001101011111101111010111101011111111010010001001001111011101101";
                    when "01101" => level_vec_out <= "1001101011111101111010111101011111111010011001001001111011101101";
                    when "01110" => level_vec_out <= "1001101011111101111010111101011111111010011001001001111011101101";
                    when "01111" => level_vec_out <= "1001101011111101111010111101011111111010011001001101111011101101";
                    when "10000" => level_vec_out <= "1001101011111101111010111101011111111010011001001101111111101101";
                    when "10001" => level_vec_out <= "1001101011111101111010111101011111111110011001001101111111101101";
                    when "10010" => level_vec_out <= "1001101011111101111010111101011111111110011001001101111111101101";
                    when "10011" => level_vec_out <= "1001101011111101111010111101011111111110011001101111111111101101";
                    when "10100" => level_vec_out <= "1001111011111101111110111101011111111110011001101111111111101101";
                    when "10101" => level_vec_out <= "1001111011111101111110111101011111111110011001101111111111101101";
                    when "10110" => level_vec_out <= "1001111011111101111110111101011111111111011001101111111111101101";
                    when "10111" => level_vec_out <= "1001111011111101111110111101011111111111011001101111111111111101";
                    when "11000" => level_vec_out <= "1001111011111111111110111101011111111111111001101111111111111101";
                    when "11001" => level_vec_out <= "1001111111111111111111111101011111111111111001101111111111111101";
                    when "11010" => level_vec_out <= "1011111111111111111111111101011111111111111001101111111111111101";
                    when "11011" => level_vec_out <= "1011111111111111111111111101011111111111111001111111111111111101";
                    when "11100" => level_vec_out <= "1011111111111111111111111101011111111111111101111111111111111111";
                    when "11101" => level_vec_out <= "1111111111111111111111111101011111111111111101111111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111101011111111111111101111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111101011111111111111101111111111111111111";
                when others => null;
                end case;
            when "010" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0001101010110101110101011110010011011100100110111000110101000011";
                    when "00001" => level_vec_out <= "0001101010110101110101011110010011011100100110111000110101000011";
                    when "00010" => level_vec_out <= "0001101010110101110101011110010011011100100110111000110101000011";
                    when "00011" => level_vec_out <= "1001101010110101110111011110010011011100100110111000110101000011";
                    when "00100" => level_vec_out <= "1001101010110101110111011110010011011100100110111000110101000011";
                    when "00101" => level_vec_out <= "1001101010110111111111011110010011011100100110111000110101000011";
                    when "00110" => level_vec_out <= "1001101010110111111111011110010011011100100110111100110101000011";
                    when "00111" => level_vec_out <= "1001101010110111111111011110010011011100100110111100110101010011";
                    when "01000" => level_vec_out <= "1001101010110111111111011110010011011100100110111101110101010011";
                    when "01001" => level_vec_out <= "1001111010110111111111011110010011011100100110111101110101010011";
                    when "01010" => level_vec_out <= "1001111010110111111111011110011011011100100110111101110101010011";
                    when "01011" => level_vec_out <= "1011111010111111111111011110011011011100100110111101110101010011";
                    when "01100" => level_vec_out <= "1011111010111111111111011110011011011100100110111101110101010011";
                    when "01101" => level_vec_out <= "1011111010111111111111011110011011011100100110111101111101010011";
                    when "01110" => level_vec_out <= "1011111010111111111111011110011011011100100110111101111101010011";
                    when "01111" => level_vec_out <= "1011111010111111111111011110011011011100100110111101111101010011";
                    when "10000" => level_vec_out <= "1011111110111111111111011110011011011100100111111101111101010011";
                    when "10001" => level_vec_out <= "1011111110111111111111011110011011011100100111111101111101110011";
                    when "10010" => level_vec_out <= "1011111110111111111111011110011011011100100111111101111101110011";
                    when "10011" => level_vec_out <= "1011111110111111111111011110011011011100100111111101111101110011";
                    when "10100" => level_vec_out <= "1011111110111111111111011110011011011100100111111101111101110011";
                    when "10101" => level_vec_out <= "1011111110111111111111011110011011011110100111111101111101110011";
                    when "10110" => level_vec_out <= "1011111110111111111111011110011011011110100111111101111101111011";
                    when "10111" => level_vec_out <= "1011111110111111111111011110011011011110100111111111111101111011";
                    when "11000" => level_vec_out <= "1011111110111111111111111110011011011110110111111111111101111011";
                    when "11001" => level_vec_out <= "1011111110111111111111111110111011011110110111111111111101111011";
                    when "11010" => level_vec_out <= "1011111110111111111111111110111011011110110111111111111111111011";
                    when "11011" => level_vec_out <= "1011111110111111111111111110111011111110111111111111111111111011";
                    when "11100" => level_vec_out <= "1011111110111111111111111110111111111110111111111111111111111011";
                    when "11101" => level_vec_out <= "1011111110111111111111111110111111111110111111111111111111111011";
                    when "11110" => level_vec_out <= "1111111110111111111111111111111111111110111111111111111111111011";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "011" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1101101010001000101111010000001010110011110000110100001101110000";
                    when "00001" => level_vec_out <= "1101101010001000101111011000001010110011110000110100001101110000";
                    when "00010" => level_vec_out <= "1101101010001000101111011000001010110011110000110110001101110000";
                    when "00011" => level_vec_out <= "1101101010001000101111011000001010110011110001110110001101110000";
                    when "00100" => level_vec_out <= "1101101011001000101111011001001010110011110001110110001101110000";
                    when "00101" => level_vec_out <= "1101101011001000101111011001001010110011110001110110001111110000";
                    when "00110" => level_vec_out <= "1101101011001000101111011001001011110011110001110110001111110000";
                    when "00111" => level_vec_out <= "1101101011001000101111011001001111111011110001110110001111110000";
                    when "01000" => level_vec_out <= "1101101011011000101111011101001111111011110011110110001111110000";
                    when "01001" => level_vec_out <= "1101101011011000101111011101011111111011110011110110001111110000";
                    when "01010" => level_vec_out <= "1101101111011000111111011101011111111011110011110110001111110000";
                    when "01011" => level_vec_out <= "1101101111011000111111011101011111111011110011110110001111110000";
                    when "01100" => level_vec_out <= "1101101111011000111111011101011111111011110011110110001111110000";
                    when "01101" => level_vec_out <= "1101101111011000111111111101011111111011110011110110001111110010";
                    when "01110" => level_vec_out <= "1101101111011001111111111101011111111111110011110110001111110010";
                    when "01111" => level_vec_out <= "1101101111011101111111111101011111111111110011110110001111110010";
                    when "10000" => level_vec_out <= "1101111111011101111111111101011111111111110011110110001111111010";
                    when "10001" => level_vec_out <= "1111111111011101111111111101011111111111110011110110001111111010";
                    when "10010" => level_vec_out <= "1111111111111111111111111101111111111111110011110110001111111010";
                    when "10011" => level_vec_out <= "1111111111111111111111111111111111111111110011110110001111111010";
                    when "10100" => level_vec_out <= "1111111111111111111111111111111111111111110011110110001111111010";
                    when "10101" => level_vec_out <= "1111111111111111111111111111111111111111111011110110011111111010";
                    when "10110" => level_vec_out <= "1111111111111111111111111111111111111111111011110110011111111111";
                    when "10111" => level_vec_out <= "1111111111111111111111111111111111111111111011110110011111111111";
                    when "11000" => level_vec_out <= "1111111111111111111111111111111111111111111111110110011111111111";
                    when "11001" => level_vec_out <= "1111111111111111111111111111111111111111111111111110011111111111";
                    when "11010" => level_vec_out <= "1111111111111111111111111111111111111111111111111110011111111111";
                    when "11011" => level_vec_out <= "1111111111111111111111111111111111111111111111111110011111111111";
                    when "11100" => level_vec_out <= "1111111111111111111111111111111111111111111111111110011111111111";
                    when "11101" => level_vec_out <= "1111111111111111111111111111111111111111111111111110111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111111111111110111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "100" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1110011111110101111100011001110100100011111110000110001101001111";
                    when "00001" => level_vec_out <= "1110011111110101111100011001110100100011111110001110001101001111";
                    when "00010" => level_vec_out <= "1110011111110101111100011001111100100011111110101110001101001111";
                    when "00011" => level_vec_out <= "1110011111110101111100011001111100100011111110101110001101001111";
                    when "00100" => level_vec_out <= "1110011111110101111100011001111100100011111110101110001101001111";
                    when "00101" => level_vec_out <= "1110011111110101111100011001111100100011111110101110011101001111";
                    when "00110" => level_vec_out <= "1110011111111101111100011001111100100011111110101110011101001111";
                    when "00111" => level_vec_out <= "1110011111111101111100011001111110100011111110101110011101001111";
                    when "01000" => level_vec_out <= "1110111111111101111100011001111110100011111110101110011101001111";
                    when "01001" => level_vec_out <= "1110111111111101111101011001111110110011111110101110011101001111";
                    when "01010" => level_vec_out <= "1110111111111101111101011001111110110011111110101111011101001111";
                    when "01011" => level_vec_out <= "1110111111111101111101011001111110110011111110101111011111001111";
                    when "01100" => level_vec_out <= "1110111111111101111101011101111110110011111110101111011111001111";
                    when "01101" => level_vec_out <= "1110111111111101111101011101111110110011111110101111011111001111";
                    when "01110" => level_vec_out <= "1110111111111101111101011101111110110011111110101111011111001111";
                    when "01111" => level_vec_out <= "1110111111111101111101011101111110110011111110101111011111001111";
                    when "10000" => level_vec_out <= "1110111111111101111101011101111110110011111110101111011111001111";
                    when "10001" => level_vec_out <= "1110111111111111111101011101111110110011111110101111011111001111";
                    when "10010" => level_vec_out <= "1110111111111111111101011101111110110011111110101111011111001111";
                    when "10011" => level_vec_out <= "1110111111111111111101011101111110110011111110101111011111001111";
                    when "10100" => level_vec_out <= "1110111111111111111101011101111110111011111110101111011111001111";
                    when "10101" => level_vec_out <= "1110111111111111111101011101111110111011111110101111011111001111";
                    when "10110" => level_vec_out <= "1110111111111111111101011101111110111011111111101111011111001111";
                    when "10111" => level_vec_out <= "1110111111111111111101011101111110111011111111101111011111101111";
                    when "11000" => level_vec_out <= "1110111111111111111101011101111110111011111111101111011111101111";
                    when "11001" => level_vec_out <= "1110111111111111111101011101111110111011111111101111011111101111";
                    when "11010" => level_vec_out <= "1110111111111111111101011111111110111011111111101111011111101111";
                    when "11011" => level_vec_out <= "1111111111111111111101011111111110111011111111101111011111101111";
                    when "11100" => level_vec_out <= "1111111111111111111111011111111110111011111111111111011111101111";
                    when "11101" => level_vec_out <= "1111111111111111111111011111111110111111111111111111011111101111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111110111111111111111111011111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111110111111111111111111111111111111";
                when others => null;
                end case;
            when "101" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1000001011010000011110011001101101000111100001100001000111101101";
                    when "00001" => level_vec_out <= "1000001011010000011110011001101101000111100001100001000111101101";
                    when "00010" => level_vec_out <= "1000101011010000011110011001101101000111100001100001000111101101";
                    when "00011" => level_vec_out <= "1000101011010000011110011001101101000111100001100001000111101101";
                    when "00100" => level_vec_out <= "1000101011010000011110011001101101000111100001100001000111101101";
                    when "00101" => level_vec_out <= "1000101011010000011110011001101101000111100001100001000111101101";
                    when "00110" => level_vec_out <= "1000101011010000011110011001101101000111100001100001000111101101";
                    when "00111" => level_vec_out <= "1000101011010000011110011001101101000111100001100001000111101101";
                    when "01000" => level_vec_out <= "1000101011010000011110011001101101000111110001100001000111101101";
                    when "01001" => level_vec_out <= "1000101011010000011110011001101101000111110001100001001111101101";
                    when "01010" => level_vec_out <= "1000101011010000011110011001101101000111110101100001001111101101";
                    when "01011" => level_vec_out <= "1000101011010000011110011001101101000111110101100001001111101101";
                    when "01100" => level_vec_out <= "1000101011010001011110011011101101000111110101100011001111101101";
                    when "01101" => level_vec_out <= "1000101011010001011110011011101101110111110101100011001111101101";
                    when "01110" => level_vec_out <= "1000101011110001111110011011101101110111110101100011001111101101";
                    when "01111" => level_vec_out <= "1100101011110001111110011011101101110111110101100111001111101101";
                    when "10000" => level_vec_out <= "1100101111110001111110011011101101110111110101100111001111101101";
                    when "10001" => level_vec_out <= "1100101111110001111110011011101101110111111101100111001111101111";
                    when "10010" => level_vec_out <= "1100101111110001111111011011101101110111111101100111011111101111";
                    when "10011" => level_vec_out <= "1100111111110001111111011011101101110111111101100111011111111111";
                    when "10100" => level_vec_out <= "1100111111110001111111011011101101110111111101110111011111111111";
                    when "10101" => level_vec_out <= "1100111111110001111111011011101101111111111101111111011111111111";
                    when "10110" => level_vec_out <= "1100111111110001111111011011101101111111111111111111011111111111";
                    when "10111" => level_vec_out <= "1100111111110101111111011011101101111111111111111111011111111111";
                    when "11000" => level_vec_out <= "1100111111110101111111011011101101111111111111111111011111111111";
                    when "11001" => level_vec_out <= "1100111111110101111111011011101101111111111111111111011111111111";
                    when "11010" => level_vec_out <= "1101111111111101111111011011101101111111111111111111011111111111";
                    when "11011" => level_vec_out <= "1101111111111111111111011111101101111111111111111111011111111111";
                    when "11100" => level_vec_out <= "1111111111111111111111011111101101111111111111111111111111111111";
                    when "11101" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "110" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0011011001110000111110101010111100100010001111111000101100010001";
                    when "00001" => level_vec_out <= "0011011001110000111110101010111100100010001111111000111100010001";
                    when "00010" => level_vec_out <= "0011011001110000111110101010111100100010001111111000111110010001";
                    when "00011" => level_vec_out <= "0011011001110000111110101010111100100010001111111000111110010001";
                    when "00100" => level_vec_out <= "1011011001110000111110101010111100100010001111111000111110010001";
                    when "00101" => level_vec_out <= "1011011001110010111110101010111100100010001111111000111110010001";
                    when "00110" => level_vec_out <= "1111011001110110111110101010111100100010001111111000111110010001";
                    when "00111" => level_vec_out <= "1111011001110110111110101010111100100010001111111000111110010001";
                    when "01000" => level_vec_out <= "1111011001110110111110101010111100100010001111111000111110010001";
                    when "01001" => level_vec_out <= "1111011001110110111110101010111100100010001111111000111110010001";
                    when "01010" => level_vec_out <= "1111011001110110111110101010111100100010001111111000111110010001";
                    when "01011" => level_vec_out <= "1111011011110110111110101010111100100010001111111000111110010101";
                    when "01100" => level_vec_out <= "1111011011110111111110101010111100100010001111111000111110010101";
                    when "01101" => level_vec_out <= "1111011011110111111110101010111100100010001111111000111110010101";
                    when "01110" => level_vec_out <= "1111011011110111111110101010111100100010001111111010111110011101";
                    when "01111" => level_vec_out <= "1111011011110111111110101010111110100010001111111010111110011101";
                    when "10000" => level_vec_out <= "1111011011110111111110101010111110100010001111111010111110111101";
                    when "10001" => level_vec_out <= "1111011111110111111110101010111110100010001111111110111110111101";
                    when "10010" => level_vec_out <= "1111011111110111111110101010111110100010001111111110111110111101";
                    when "10011" => level_vec_out <= "1111011111110111111110101010111110110010001111111110111110111101";
                    when "10100" => level_vec_out <= "1111011111111111111110101010111111110010001111111110111110111111";
                    when "10101" => level_vec_out <= "1111011111111111111110101010111111110010011111111110111110111111";
                    when "10110" => level_vec_out <= "1111011111111111111110101010111111110010011111111111111110111111";
                    when "10111" => level_vec_out <= "1111011111111111111110101010111111110010011111111111111110111111";
                    when "11000" => level_vec_out <= "1111011111111111111110101010111111110010111111111111111110111111";
                    when "11001" => level_vec_out <= "1111111111111111111110101010111111110010111111111111111110111111";
                    when "11010" => level_vec_out <= "1111111111111111111110111011111111110010111111111111111110111111";
                    when "11011" => level_vec_out <= "1111111111111111111110111011111111110110111111111111111111111111";
                    when "11100" => level_vec_out <= "1111111111111111111110111011111111110110111111111111111111111111";
                    when "11101" => level_vec_out <= "1111111111111111111110111011111111110110111111111111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111110111011111111110111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111011111111111111111111111111111111111111";
                when others => null;
                end case;
            when "111" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1010101000111001011010110100000011011100001100111000001001100011";
                    when "00001" => level_vec_out <= "1010101000111001011010110100000011011100001111111000001001100011";
                    when "00010" => level_vec_out <= "1010101000111001111010110100000011011100001111111010001001100011";
                    when "00011" => level_vec_out <= "1010101000111001111010110110000011011100001111111010001001100011";
                    when "00100" => level_vec_out <= "1010101000111001111010110110000111011100001111111010001001100011";
                    when "00101" => level_vec_out <= "1010101000111001111010110110000111011100001111111010001001100011";
                    when "00110" => level_vec_out <= "1010101000111001111010110110000111011110001111111010001001100011";
                    when "00111" => level_vec_out <= "1010101000111101111010110110000111011110001111111010001001100011";
                    when "01000" => level_vec_out <= "1010111000111101111010110110000111011110001111111010001001100011";
                    when "01001" => level_vec_out <= "1010111000111101111010110110000111011110011111111010001001100011";
                    when "01010" => level_vec_out <= "1010111100111101111010110110100111011110011111111110001001100011";
                    when "01011" => level_vec_out <= "1010111100111101111110110110100111011110011111111110001001100111";
                    when "01100" => level_vec_out <= "1010111100111101111110110110100111011110011111111110001001100111";
                    when "01101" => level_vec_out <= "1010111100111101111110110110101111011110011111111110101001100111";
                    when "01110" => level_vec_out <= "1110111100111101111110110110101111011110011111111110101001100111";
                    when "01111" => level_vec_out <= "1110111100111101111110110110111111011111011111111110111001100111";
                    when "10000" => level_vec_out <= "1110111100111101111110110110111111011111011111111110111001100111";
                    when "10001" => level_vec_out <= "1110111100111101111110110110111111011111011111111110111001100111";
                    when "10010" => level_vec_out <= "1110111100111111111110110110111111011111011111111110111001111111";
                    when "10011" => level_vec_out <= "1110111100111111111110110110111111011111011111111110111001111111";
                    when "10100" => level_vec_out <= "1110111100111111111110110110111111011111011111111110111011111111";
                    when "10101" => level_vec_out <= "1110111101111111111110110110111111011111011111111110111011111111";
                    when "10110" => level_vec_out <= "1110111101111111111110110110111111011111111111111110111011111111";
                    when "10111" => level_vec_out <= "1111111111111111111110111111111111011111111111111110111011111111";
                    when "11000" => level_vec_out <= "1111111111111111111110111111111111011111111111111111111011111111";
                    when "11001" => level_vec_out <= "1111111111111111111110111111111111011111111111111111111011111111";
                    when "11010" => level_vec_out <= "1111111111111111111110111111111111111111111111111111111011111111";
                    when "11011" => level_vec_out <= "1111111111111111111110111111111111111111111111111111111011111111";
                    when "11100" => level_vec_out <= "1111111111111111111110111111111111111111111111111111111011111111";
                    when "11101" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111011111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111011111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111011111111";
                when others => null;
                end case;
            when others => null;
        end case;
    end process;
end Behavioral;