/**
 * @file level_hvec_gen_hdl.hpp
 * @brief This script generates HDL code for generating high-dimensional LEVEL vectors.
 * It is a novel method; for more information, please refer to our paper.
 *
 * @author Saeid Jamili and Marco Angioli
 * @note Author names are listed in alphabetical order.
 * @email <saeid.jamili@uniroma1.it>
 * @email <marco.angioli@uniroma1.it>
 *
 * @contributors
 *
 * @date Created: 24th July 2023
 * @date Last Updated: 23th August 2023
 *
 * @version 1.0.0
 *
 * @institute Sapienza University of Rome
 * @cite https://doi.org/10.xxxx/yyyyy
 *
 * @section DEPENDENCIES
 * - Dependency1: Description or version details.
 * - Dependency2: Description or version details.
 *
 * @section LICENSE
 * This file is part of the Aeneas HyperCompute Platform.
 *
 * Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 *
 * @section CHANGELOG
 * @version 1.0.0-dev - 23th August 2023
 * - Initial release
 *
 * @todo
 * - Complete level vector generator function
 * - Add training
 *
 * @see
 * -
 * -
 * -
 *
 */

module level_vec_gen (
    output reg [63:0] level_vec_out,
    input [2:0] frame_index,
    input [4:0] frame_id
);
    always @(*) begin
        // Update this function to match your requirements
        case (frame_index)
            0: begin
                case (frame_id)
                    0: level_vec_out = 64'b1100100101000110000111011100101011100001111000000111010110000110;
                    1: level_vec_out = 64'b1100100101000110010111011100101011100001111000000111010110001110;
                    2: level_vec_out = 64'b1100100101000110011111011100101011100001111010000111011110001110;
                    3: level_vec_out = 64'b1100100101000110011111011100101011100001111011000111011110001110;
                    4: level_vec_out = 64'b1100100101000110011111011100101011100001111011000111011110001110;
                    5: level_vec_out = 64'b1110100101000110011111011100101011100001111011000111011110001110;
                    6: level_vec_out = 64'b1110100101000110011111011100101011100001111011000111011110001110;
                    7: level_vec_out = 64'b1110100101000110011111111100101011100001111011000111011110001110;
                    8: level_vec_out = 64'b1110100101000110011111111100101111100001111011000111011110001110;
                    9: level_vec_out = 64'b1110100101000110011111111100101111100001111011000111011110001110;
                    10: level_vec_out = 64'b1110100101000110011111111100101111110001111011000111011110001110;
                    11: level_vec_out = 64'b1110100101000110011111111100101111110001111011000111011110001110;
                    12: level_vec_out = 64'b1110100101000110011111111100101111110001111011010111011110011110;
                    13: level_vec_out = 64'b1110100111000110111111111100101111111001111011010111011110011110;
                    14: level_vec_out = 64'b1110101111000110111111111100101111111001111011110111011110011110;
                    15: level_vec_out = 64'b1110101111000110111111111100101111111001111011111111011110111110;
                    16: level_vec_out = 64'b1110101111010110111111111100101111111001111011111111011110111110;
                    17: level_vec_out = 64'b1110101111110110111111111100101111111001111011111111011110111110;
                    18: level_vec_out = 64'b1110101111110110111111111100101111111001111011111111011110111110;
                    19: level_vec_out = 64'b1110101111110110111111111100101111111001111011111111011110111110;
                    20: level_vec_out = 64'b1110101111110110111111111100101111111011111011111111011110111110;
                    21: level_vec_out = 64'b1110101111110110111111111100101111111011111011111111011111111111;
                    22: level_vec_out = 64'b1110101111110110111111111100101111111011111111111111011111111111;
                    23: level_vec_out = 64'b1110111111110110111111111100101111111011111111111111011111111111;
                    24: level_vec_out = 64'b1110111111110110111111111110111111111011111111111111011111111111;
                    25: level_vec_out = 64'b1110111111110110111111111110111111111011111111111111011111111111;
                    26: level_vec_out = 64'b1110111111110110111111111110111111111011111111111111011111111111;
                    27: level_vec_out = 64'b1110111111110110111111111111111111111011111111111111011111111111;
                    28: level_vec_out = 64'b1110111111110110111111111111111111111011111111111111011111111111;
                    29: level_vec_out = 64'b1110111111110110111111111111111111111011111111111111011111111111;
                    30: level_vec_out = 64'b1111111111111110111111111111111111111011111111111111011111111111;
                    31: level_vec_out = 64'b1111111111111110111111111111111111111011111111111111011111111111;
                endcase
            end
            1: begin
                case (frame_id)
                    0: level_vec_out = 64'b0011011100100010111101010110001011001111100110110101000111010010;
                    1: level_vec_out = 64'b0011011100100010111101010110001011001111100110110101000111010010;
                    2: level_vec_out = 64'b0011011100100010111101010110001011001111100110110101000111010010;
                    3: level_vec_out = 64'b0011011100100011111101010111001011001111101110110101001111010010;
                    4: level_vec_out = 64'b0011011100100011111101010111001011001111101110110101001111010010;
                    5: level_vec_out = 64'b0011011100100011111101010111001011001111101110110101001111010010;
                    6: level_vec_out = 64'b0011011100100011111101010111001011001111101110110101101111010010;
                    7: level_vec_out = 64'b0011011100100011111101010111001011001111101110110101101111010010;
                    8: level_vec_out = 64'b0011011100100011111101110111001011001111101111110101101111010110;
                    9: level_vec_out = 64'b0011011100100011111101110111001011001111101111110101101111010110;
                    10: level_vec_out = 64'b0011011100100011111101110111011011001111101111110101101111010110;
                    11: level_vec_out = 64'b0011011100100011111101111111011111001111101111110101101111010110;
                    12: level_vec_out = 64'b0011111100100011111101111111011111001111101111111101101111010110;
                    13: level_vec_out = 64'b0011111100100011111101111111011111001111101111111101101111010110;
                    14: level_vec_out = 64'b0011111100100011111101111111011111001111101111111101101111110110;
                    15: level_vec_out = 64'b0011111100110011111101111111011111011111101111111101101111110110;
                    16: level_vec_out = 64'b0011111100110011111101111111111111011111101111111101101111110110;
                    17: level_vec_out = 64'b0011111100110011111101111111111111011111101111111101101111110110;
                    18: level_vec_out = 64'b0011111100110011111101111111111111011111101111111101101111110110;
                    19: level_vec_out = 64'b0011111110110011111101111111111111011111101111111101101111110110;
                    20: level_vec_out = 64'b0011111110110011111101111111111111011111101111111101101111110110;
                    21: level_vec_out = 64'b0011111110110011111111111111111111011111101111111101101111110111;
                    22: level_vec_out = 64'b0011111110110011111111111111111111011111101111111111101111110111;
                    23: level_vec_out = 64'b0011111110111011111111111111111111011111101111111111101111110111;
                    24: level_vec_out = 64'b0011111110111011111111111111111111011111101111111111101111110111;
                    25: level_vec_out = 64'b0111111110111011111111111111111111011111111111111111101111110111;
                    26: level_vec_out = 64'b1111111111111011111111111111111111011111111111111111101111111111;
                    27: level_vec_out = 64'b1111111111111011111111111111111111011111111111111111111111111111;
                    28: level_vec_out = 64'b1111111111111011111111111111111111011111111111111111111111111111;
                    29: level_vec_out = 64'b1111111111111011111111111111111111111111111111111111111111111111;
                    30: level_vec_out = 64'b1111111111111011111111111111111111111111111111111111111111111111;
                    31: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                endcase
            end
            2: begin
                case (frame_id)
                    0: level_vec_out = 64'b1100110111001010101100110100000001111010001011110101011110000110;
                    1: level_vec_out = 64'b1100110111001010101110110100000001111010001011110101011110000110;
                    2: level_vec_out = 64'b1100110111001010101110110100000001111010001011110101011110000110;
                    3: level_vec_out = 64'b1100110111001010101110110100000011111010001011110101011110000110;
                    4: level_vec_out = 64'b1100110111011010101110110110000011111010001011110101011110000110;
                    5: level_vec_out = 64'b1100110111011010101110110110000011111110001011110101011110000110;
                    6: level_vec_out = 64'b1100110111011010111110110110000011111110001011110101011110010110;
                    7: level_vec_out = 64'b1100111111011010111110110110000011111110001011110101011110010110;
                    8: level_vec_out = 64'b1100111111011010111111110110000011111110001011110101011110010110;
                    9: level_vec_out = 64'b1100111111011010111111110110000011111110101011110101011110010110;
                    10: level_vec_out = 64'b1100111111011010111111110110000011111110101011110101011110010110;
                    11: level_vec_out = 64'b1100111111111010111111110110000011111110101011110101111110010110;
                    12: level_vec_out = 64'b1100111111111010111111110110000011111110101011110101111110010110;
                    13: level_vec_out = 64'b1100111111111010111111110110010011111111101111110101111110010110;
                    14: level_vec_out = 64'b1110111111111010111111110110010011111111101111110101111110010110;
                    15: level_vec_out = 64'b1110111111111010111111110110010011111111101111110101111110010110;
                    16: level_vec_out = 64'b1110111111111010111111111110010011111111111111110101111110010110;
                    17: level_vec_out = 64'b1111111111111011111111111110010011111111111111110101111110011110;
                    18: level_vec_out = 64'b1111111111111011111111111110010011111111111111110101111110011110;
                    19: level_vec_out = 64'b1111111111111011111111111111010011111111111111110101111110011110;
                    20: level_vec_out = 64'b1111111111111011111111111111110011111111111111110101111110011110;
                    21: level_vec_out = 64'b1111111111111011111111111111110011111111111111110101111110011110;
                    22: level_vec_out = 64'b1111111111111011111111111111110011111111111111110101111110011110;
                    23: level_vec_out = 64'b1111111111111011111111111111110111111111111111110101111111011110;
                    24: level_vec_out = 64'b1111111111111011111111111111110111111111111111110101111111011110;
                    25: level_vec_out = 64'b1111111111111011111111111111110111111111111111110111111111011110;
                    26: level_vec_out = 64'b1111111111111011111111111111110111111111111111110111111111011111;
                    27: level_vec_out = 64'b1111111111111011111111111111110111111111111111110111111111111111;
                    28: level_vec_out = 64'b1111111111111011111111111111110111111111111111111111111111111111;
                    29: level_vec_out = 64'b1111111111111011111111111111110111111111111111111111111111111111;
                    30: level_vec_out = 64'b1111111111111011111111111111110111111111111111111111111111111111;
                    31: level_vec_out = 64'b1111111111111011111111111111110111111111111111111111111111111111;
                endcase
            end
            3: begin
                case (frame_id)
                    0: level_vec_out = 64'b0010001000100101011111100010100010001010101001110100111010110100;
                    1: level_vec_out = 64'b0011001000100101111111100010100010001010101001110100111010110100;
                    2: level_vec_out = 64'b0011001000100101111111100010100010001010101001110100111010110100;
                    3: level_vec_out = 64'b0011001000100101111111100010100010001010101001110100111010110100;
                    4: level_vec_out = 64'b0011001000100101111111100010100110001010101011110100111010110100;
                    5: level_vec_out = 64'b0011001000100101111111100010100110001010101011110100111010110100;
                    6: level_vec_out = 64'b0011011000100101111111100010100110001010101011110100111010110100;
                    7: level_vec_out = 64'b0011011000100111111111100010100110001010101011110100111010110100;
                    8: level_vec_out = 64'b0011011001101111111111100010100110001010101011110100111010110100;
                    9: level_vec_out = 64'b0011011001101111111111100010100110001010101011111100111010110100;
                    10: level_vec_out = 64'b0011011001101111111111100010100110001010101011111100111110110100;
                    11: level_vec_out = 64'b0011011001101111111111100010100110001010101011111100111110110100;
                    12: level_vec_out = 64'b0011011001101111111111100010100110001010101011111100111110110100;
                    13: level_vec_out = 64'b0011011001101111111111100010100110001010101011111100111110110100;
                    14: level_vec_out = 64'b0011011001101111111111100010100110001010111011111100111110110100;
                    15: level_vec_out = 64'b0011011001101111111111100010100110001010111011111100111110110100;
                    16: level_vec_out = 64'b1011011001101111111111100110100110001010111011111100111110110100;
                    17: level_vec_out = 64'b1011011001101111111111100110100110001010111011111100111110110100;
                    18: level_vec_out = 64'b1011011001101111111111110110110110001010111011111100111110111100;
                    19: level_vec_out = 64'b1011011001101111111111110111110110001010111011111100111110111100;
                    20: level_vec_out = 64'b1011011001101111111111110111110110101010111011111100111111111110;
                    21: level_vec_out = 64'b1011011101101111111111110111110110101010111011111100111111111110;
                    22: level_vec_out = 64'b1011111101101111111111110111110110101010111011111100111111111111;
                    23: level_vec_out = 64'b1011111101101111111111110111110110101010111011111100111111111111;
                    24: level_vec_out = 64'b1011111111101111111111111111110110101010111011111100111111111111;
                    25: level_vec_out = 64'b1011111111101111111111111111110110101010111111111100111111111111;
                    26: level_vec_out = 64'b1111111111101111111111111111110110101010111111111100111111111111;
                    27: level_vec_out = 64'b1111111111101111111111111111110110111110111111111100111111111111;
                    28: level_vec_out = 64'b1111111111101111111111111111110110111110111111111100111111111111;
                    29: level_vec_out = 64'b1111111111101111111111111111110110111110111111111101111111111111;
                    30: level_vec_out = 64'b1111111111111111111111111111110111111110111111111101111111111111;
                    31: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                endcase
            end
            4: begin
                case (frame_id)
                    0: level_vec_out = 64'b0011010000100011101101010010010100111100111000101101110100011010;
                    1: level_vec_out = 64'b0011010000100011101101010010011100111100111000101101110100011010;
                    2: level_vec_out = 64'b1011010000100011101101010010011100111100111000111101110100011010;
                    3: level_vec_out = 64'b1011010000100011101101010010011100111100111000111101110100011010;
                    4: level_vec_out = 64'b1011010000100011101101010010011100111100111000111101110100011011;
                    5: level_vec_out = 64'b1011010001100011101101010010011110111100111000111101110100011011;
                    6: level_vec_out = 64'b1011010001100011101101010010011110111100111000111101110100011011;
                    7: level_vec_out = 64'b1111010001110011101101010010011110111100111000111101110100011011;
                    8: level_vec_out = 64'b1111010001110011101101010010011110111100111000111101110100011011;
                    9: level_vec_out = 64'b1111010011110011101101010010011110111100111001111101110100011011;
                    10: level_vec_out = 64'b1111010011110011101101010010011110111100111001111101110100011011;
                    11: level_vec_out = 64'b1111010011110011101101010010011110111100111001111101110100011011;
                    12: level_vec_out = 64'b1111010011110011101101011010011111111100111001111101110100011011;
                    13: level_vec_out = 64'b1111010011111011101101011010011111111100111001111101110100011011;
                    14: level_vec_out = 64'b1111010011111011101101011010011111111100111001111101110100011011;
                    15: level_vec_out = 64'b1111011011111011101101011011011111111100111001111101110101011011;
                    16: level_vec_out = 64'b1111011011111011101101011011011111111100111001111101110101111011;
                    17: level_vec_out = 64'b1111111011111011101101011011011111111100111001111101110101111011;
                    18: level_vec_out = 64'b1111111011111011101101011011011111111100111001111101110101111011;
                    19: level_vec_out = 64'b1111111011111011101101011011011111111110111101111101110101111011;
                    20: level_vec_out = 64'b1111111011111011101101011011011111111110111101111101110101111011;
                    21: level_vec_out = 64'b1111111011111011101101011011011111111110111101111101110101111011;
                    22: level_vec_out = 64'b1111111111111011101101011011011111111110111101111101110111111011;
                    23: level_vec_out = 64'b1111111111111011101101011011011111111110111101111111110111111111;
                    24: level_vec_out = 64'b1111111111111011101101011111011111111110111101111111110111111111;
                    25: level_vec_out = 64'b1111111111111011101101011111011111111111111111111111110111111111;
                    26: level_vec_out = 64'b1111111111111011111111011111011111111111111111111111110111111111;
                    27: level_vec_out = 64'b1111111111111011111111011111011111111111111111111111110111111111;
                    28: level_vec_out = 64'b1111111111111011111111011111111111111111111111111111110111111111;
                    29: level_vec_out = 64'b1111111111111111111111011111111111111111111111111111110111111111;
                    30: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    31: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                endcase
            end
            5: begin
                case (frame_id)
                    0: level_vec_out = 64'b0011101111100001110001010100000100001110100001011011101001101011;
                    1: level_vec_out = 64'b0011101111100001110001011100000100001110100001011011101001101011;
                    2: level_vec_out = 64'b0011101111100001110001011100000100001110100001111011101001101011;
                    3: level_vec_out = 64'b0011111111100001110001011100000100001110100001111011101001101011;
                    4: level_vec_out = 64'b0011111111100001110001011100000100001110100001111011101001101011;
                    5: level_vec_out = 64'b0011111111100001110001011100000100001110100001111011101001101011;
                    6: level_vec_out = 64'b0011111111100101110001011100001100001111100001111011101001101011;
                    7: level_vec_out = 64'b0011111111100101110001011100001100011111100001111011101001101011;
                    8: level_vec_out = 64'b0011111111100101110001011100001100011111100001111011101001101011;
                    9: level_vec_out = 64'b0011111111100101110001011100101100011111100001111011101001101011;
                    10: level_vec_out = 64'b0011111111100101110001011100101101011111100001111111111001101011;
                    11: level_vec_out = 64'b0011111111100101110001011100101111011111100001111111111001101011;
                    12: level_vec_out = 64'b0011111111100101110001011100101111011111100001111111111001101011;
                    13: level_vec_out = 64'b0011111111100101110001011100101111011111100001111111111001101011;
                    14: level_vec_out = 64'b0011111111100101110001011100111111011111100001111111111001101011;
                    15: level_vec_out = 64'b0011111111100101110001011100111111011111100001111111111001101011;
                    16: level_vec_out = 64'b0011111111100101110001011100111111011111100001111111111001101011;
                    17: level_vec_out = 64'b0011111111100101110001111100111111011111100001111111111001101011;
                    18: level_vec_out = 64'b0111111111101101110101111100111111011111100001111111111001101011;
                    19: level_vec_out = 64'b0111111111101101110101111100111111011111100001111111111001101111;
                    20: level_vec_out = 64'b0111111111101101110101111110111111011111110001111111111001101111;
                    21: level_vec_out = 64'b0111111111101101111111111110111111011111110001111111111001101111;
                    22: level_vec_out = 64'b1111111111101101111111111110111111011111110001111111111001101111;
                    23: level_vec_out = 64'b1111111111101101111111111111111111011111110001111111111001101111;
                    24: level_vec_out = 64'b1111111111101101111111111111111111011111110001111111111001101111;
                    25: level_vec_out = 64'b1111111111101101111111111111111111011111110001111111111001101111;
                    26: level_vec_out = 64'b1111111111101101111111111111111111011111110001111111111001101111;
                    27: level_vec_out = 64'b1111111111101101111111111111111111111111110001111111111001101111;
                    28: level_vec_out = 64'b1111111111111101111111111111111111111111110101111111111111101111;
                    29: level_vec_out = 64'b1111111111111101111111111111111111111111111111111111111111101111;
                    30: level_vec_out = 64'b1111111111111101111111111111111111111111111111111111111111101111;
                    31: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111101111;
                endcase
            end
            6: begin
                case (frame_id)
                    0: level_vec_out = 64'b1100101000110110111101100010000110110110001001011001011111100111;
                    1: level_vec_out = 64'b1100101000110110111101100010000110110110001001011001011111100111;
                    2: level_vec_out = 64'b1100101000111110111101100010000110110110001001011001011111100111;
                    3: level_vec_out = 64'b1100101000111110111101100010000110110110001001011001011111100111;
                    4: level_vec_out = 64'b1100101000111110111101110010000110110110001001011011011111100111;
                    5: level_vec_out = 64'b1100101000111110111101110110000110110110001001011011011111100111;
                    6: level_vec_out = 64'b1100101000111111111101110110000110110110001001011011011111100111;
                    7: level_vec_out = 64'b1100101000111111111101110110000110110110011001011011011111100111;
                    8: level_vec_out = 64'b1100101000111111111101110110000110110110011001011011011111100111;
                    9: level_vec_out = 64'b1100101010111111111101110110000110110110011001011011011111101111;
                    10: level_vec_out = 64'b1100101010111111111101110111000110110110011001011011011111101111;
                    11: level_vec_out = 64'b1100101010111111111101110111000111110110011001011011011111101111;
                    12: level_vec_out = 64'b1100101010111111111101111111000111110110011001011011011111101111;
                    13: level_vec_out = 64'b1100101010111111111101111111000111111110011001011011011111101111;
                    14: level_vec_out = 64'b1100101010111111111101111111000111111110011001111011011111101111;
                    15: level_vec_out = 64'b1100101010111111111101111111000111111110011001111011011111101111;
                    16: level_vec_out = 64'b1100101010111111111101111111000111111110011001111011011111101111;
                    17: level_vec_out = 64'b1100101010111111111101111111000111111110011001111011111111101111;
                    18: level_vec_out = 64'b1100101110111111111101111111000111111110011101111011111111101111;
                    19: level_vec_out = 64'b1100101110111111111101111111001111111110011101111011111111101111;
                    20: level_vec_out = 64'b1100101110111111111101111111011111111110011101111011111111101111;
                    21: level_vec_out = 64'b1100101110111111111101111111011111111110011101111011111111101111;
                    22: level_vec_out = 64'b1100101111111111111101111111011111111110011101111011111111101111;
                    23: level_vec_out = 64'b1100101111111111111101111111011111111110011101111011111111101111;
                    24: level_vec_out = 64'b1100111111111111111101111111111111111111011101111011111111101111;
                    25: level_vec_out = 64'b1100111111111111111101111111111111111111011101111011111111101111;
                    26: level_vec_out = 64'b1100111111111111111101111111111111111111011101111011111111101111;
                    27: level_vec_out = 64'b1100111111111111111101111111111111111111011101111011111111101111;
                    28: level_vec_out = 64'b1100111111111111111101111111111111111111011101111111111111101111;
                    29: level_vec_out = 64'b1110111111111111111101111111111111111111111101111111111111111111;
                    30: level_vec_out = 64'b1110111111111111111111111111111111111111111101111111111111111111;
                    31: level_vec_out = 64'b1110111111111111111111111111111111111111111101111111111111111111;
                endcase
            end
            7: begin
                case (frame_id)
                    0: level_vec_out = 64'b0111000110011011100100011111011111010110100110010110000110000001;
                    1: level_vec_out = 64'b0111000110011011100110011111011111010110100110010110000110000001;
                    2: level_vec_out = 64'b0111000110011011100110011111011111010111100110010110000110000001;
                    3: level_vec_out = 64'b0111000110011011100110011111111111010111100110010110000110000001;
                    4: level_vec_out = 64'b0111000110011011100110011111111111010111100110010110000110000011;
                    5: level_vec_out = 64'b0111100110111011100111011111111111010111100110010110000110000011;
                    6: level_vec_out = 64'b0111100110111011100111011111111111010111100110010110000110000011;
                    7: level_vec_out = 64'b0111100110111011100111111111111111010111100110010110000110000011;
                    8: level_vec_out = 64'b0111100110111011100111111111111111011111100110010110000110000011;
                    9: level_vec_out = 64'b0111100110111011100111111111111111011111100110010110000110000111;
                    10: level_vec_out = 64'b0111100110111011100111111111111111111111100110010110000110000111;
                    11: level_vec_out = 64'b0111110110111011100111111111111111111111110110010110000110000111;
                    12: level_vec_out = 64'b0111111110111011100111111111111111111111110110010110000110000111;
                    13: level_vec_out = 64'b0111111110111011100111111111111111111111110110010110000110000111;
                    14: level_vec_out = 64'b0111111110111011100111111111111111111111110110110110000110000111;
                    15: level_vec_out = 64'b0111111110111011100111111111111111111111110110110110010110000111;
                    16: level_vec_out = 64'b1111111110111011100111111111111111111111110110110110010110000111;
                    17: level_vec_out = 64'b1111111110111011101111111111111111111111110110110110010110000111;
                    18: level_vec_out = 64'b1111111110111011101111111111111111111111110110110110010110000111;
                    19: level_vec_out = 64'b1111111110111011111111111111111111111111110110110110010110000111;
                    20: level_vec_out = 64'b1111111110111011111111111111111111111111110110110110010110000111;
                    21: level_vec_out = 64'b1111111110111011111111111111111111111111110110110110110110000111;
                    22: level_vec_out = 64'b1111111110111011111111111111111111111111110110110110110110000111;
                    23: level_vec_out = 64'b1111111110111011111111111111111111111111110110110110110111000111;
                    24: level_vec_out = 64'b1111111110111011111111111111111111111111110110110110110111000111;
                    25: level_vec_out = 64'b1111111111111011111111111111111111111111110110111110110111000111;
                    26: level_vec_out = 64'b1111111111111011111111111111111111111111110110111111110111000111;
                    27: level_vec_out = 64'b1111111111111011111111111111111111111111110110111111110111011111;
                    28: level_vec_out = 64'b1111111111111011111111111111111111111111110110111111111111011111;
                    29: level_vec_out = 64'b1111111111111011111111111111111111111111110110111111111111011111;
                    30: level_vec_out = 64'b1111111111111111111111111111111111111111110110111111111111011111;
                    31: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                endcase
            end
        endcase
    end
endmodule