/**
 * @file level_hvec_gen_hdl.hpp
 * @brief This script generates HDL code for generating high-dimensional LEVEL vectors.
 * It is a novel method; for more information, please refer to our paper.
 *
 * @author Saeid Jamili and Marco Angioli
 * @note Author names are listed in alphabetical order.
 * @email <saeid.jamili@uniroma1.it>
 * @email <marco.angioli@uniroma1.it>
 *
 * @contributors
 *
 * @date Created: 24th July 2023
 * @date Last Updated: 23th August 2023
 *
 * @version 1.0.0
 *
 * @institute Sapienza University of Rome
 * @cite https://doi.org/10.xxxx/yyyyy
 *
 * @section DEPENDENCIES
 * - Dependency1: Description or version details.
 * - Dependency2: Description or version details.
 *
 * @section LICENSE
 * This file is part of the Aeneas HyperCompute Platform.
 *
 * Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 *
 * @section CHANGELOG
 * @version 1.0.0-dev - 23th August 2023
 * - Initial release
 *
 * @todo
 * - Complete level vector generator function
 * - Add training
 *
 * @see
 * -
 * -
 * -
 *
 */

module level_vec_gen (
    output reg [63:0] level_vec_out,
    input [2:0] frame_index,
    input [4:0] frame_id
);
    always @(*) begin
        // Update this function to match your requirements
        case (frame_index)
            0: begin
                case (frame_id)
                    0: level_vec_out = 64'b1111110101000000111110100100110111110100110000111000110010000011;
                    1: level_vec_out = 64'b1111110101000000111110100100110111110100110000111000110010000011;
                    2: level_vec_out = 64'b1111110101000100111110100110110111110100110000111000110010000011;
                    3: level_vec_out = 64'b1111110101010100111110100110110111111100110000111000110010000011;
                    4: level_vec_out = 64'b1111110101010100111110100110110111111100110000111001110010010011;
                    5: level_vec_out = 64'b1111110101010101111110100110110111111100110000111001110010010011;
                    6: level_vec_out = 64'b1111110101010101111110100110110111111100110000111001111010010011;
                    7: level_vec_out = 64'b1111110101110101111110100110110111111100110000111001111010010011;
                    8: level_vec_out = 64'b1111110101110101111110100110110111111100110000111001111010010111;
                    9: level_vec_out = 64'b1111110101110101111110100110110111111100110000111001111010010111;
                    10: level_vec_out = 64'b1111110101110101111110100110110111111100110000111001111010010111;
                    11: level_vec_out = 64'b1111110101110101111110100110110111111100110000111001111110011111;
                    12: level_vec_out = 64'b1111110101111101111110100110110111111100110000111001111110011111;
                    13: level_vec_out = 64'b1111110101111101111110100110110111111100110000111001111110011111;
                    14: level_vec_out = 64'b1111110101111101111110100110110111111101110010111001111110011111;
                    15: level_vec_out = 64'b1111110101111101111110110110110111111101110010111001111110011111;
                    16: level_vec_out = 64'b1111110101111101111110110110110111111111110010111001111110011111;
                    17: level_vec_out = 64'b1111110101111101111110111110110111111111110010111001111110011111;
                    18: level_vec_out = 64'b1111111101111101111110111110110111111111110010111101111110011111;
                    19: level_vec_out = 64'b1111111101111101111110111110110111111111110010111101111110111111;
                    20: level_vec_out = 64'b1111111101111101111110111110110111111111110010111101111110111111;
                    21: level_vec_out = 64'b1111111101111101111110111110110111111111110010111101111110111111;
                    22: level_vec_out = 64'b1111111101111101111110111110110111111111110011111101111110111111;
                    23: level_vec_out = 64'b1111111101111111111110111110110111111111110011111101111110111111;
                    24: level_vec_out = 64'b1111111101111111111110111110110111111111111011111101111110111111;
                    25: level_vec_out = 64'b1111111111111111111111111110110111111111111011111101111110111111;
                    26: level_vec_out = 64'b1111111111111111111111111110110111111111111011111101111110111111;
                    27: level_vec_out = 64'b1111111111111111111111111110110111111111111011111101111111111111;
                    28: level_vec_out = 64'b1111111111111111111111111110111111111111111011111101111111111111;
                    29: level_vec_out = 64'b1111111111111111111111111110111111111111111011111101111111111111;
                    30: level_vec_out = 64'b1111111111111111111111111111111111111111111011111111111111111111;
                    31: level_vec_out = 64'b1111111111111111111111111111111111111111111011111111111111111111;
                endcase
            end
            1: begin
                case (frame_id)
                    0: level_vec_out = 64'b0111001001101101110000011010100100010001111110000100100011011010;
                    1: level_vec_out = 64'b0111001001101101110100011010101100010001111110000100100011011010;
                    2: level_vec_out = 64'b0111001001101101110100011010101100010001111110000100100011011011;
                    3: level_vec_out = 64'b0111001001101101110100011010101100010001111110000100100011011011;
                    4: level_vec_out = 64'b0111001001101101110100011010101100010001111110000100100011011011;
                    5: level_vec_out = 64'b0111001001101101110100011010101100011001111110000100100011111011;
                    6: level_vec_out = 64'b0111001001101101110100011010101100011001111110000100100011111011;
                    7: level_vec_out = 64'b0111001001101101110100011010101100011001111110000100100011111011;
                    8: level_vec_out = 64'b0111101001101101110100011010101100011001111110000100111011111011;
                    9: level_vec_out = 64'b0111101001101101110100011010101100011001111110000100111011111011;
                    10: level_vec_out = 64'b0111101001101111110100011111101100011001111110000100111011111011;
                    11: level_vec_out = 64'b0111101001101111110100011111101100011001111110000100111011111011;
                    12: level_vec_out = 64'b0111101001101111110100011111101110011001111110000100111011111011;
                    13: level_vec_out = 64'b0111101001101111111100011111101110011001111110110100111011111011;
                    14: level_vec_out = 64'b0111111001101111111100011111101110011001111111110100111011111011;
                    15: level_vec_out = 64'b0111111001101111111100011111101110011001111111110100111011111011;
                    16: level_vec_out = 64'b0111111001101111111100011111101110011001111111110110111011111011;
                    17: level_vec_out = 64'b0111111001101111111100011111101110011001111111110110111011111011;
                    18: level_vec_out = 64'b0111111001101111111100011111101110011001111111110110111011111111;
                    19: level_vec_out = 64'b0111111001101111111100011111101110011011111111110110111011111111;
                    20: level_vec_out = 64'b0111111001101111111100011111101111011011111111110111111011111111;
                    21: level_vec_out = 64'b0111111101101111111100011111101111011111111111110111111011111111;
                    22: level_vec_out = 64'b0111111101101111111100011111101111011111111111110111111011111111;
                    23: level_vec_out = 64'b0111111111101111111100011111101111011111111111110111111011111111;
                    24: level_vec_out = 64'b0111111111101111111100011111101111011111111111111111111011111111;
                    25: level_vec_out = 64'b0111111111101111111110011111101111011111111111111111111011111111;
                    26: level_vec_out = 64'b0111111111101111111110011111111111011111111111111111111011111111;
                    27: level_vec_out = 64'b0111111111101111111111011111111111011111111111111111111011111111;
                    28: level_vec_out = 64'b0111111111101111111111011111111111011111111111111111111011111111;
                    29: level_vec_out = 64'b0111111111101111111111111111111111011111111111111111111011111111;
                    30: level_vec_out = 64'b0111111111111111111111111111111111111111111111111111111011111111;
                    31: level_vec_out = 64'b0111111111111111111111111111111111111111111111111111111111111111;
                endcase
            end
            2: begin
                case (frame_id)
                    0: level_vec_out = 64'b0011111000111100011010100100011110101110110100001000000100001000;
                    1: level_vec_out = 64'b0011111000111100011010100100011110101110110100001000000100001100;
                    2: level_vec_out = 64'b1011111000111100011010100100011110101110110100001000000100001101;
                    3: level_vec_out = 64'b1011111000111100011010100100011110101110110100001001000100001101;
                    4: level_vec_out = 64'b1011111000111100011010100100011110101110110100001001000100001101;
                    5: level_vec_out = 64'b1011111000111110011010100100011110101110110100001001000100101101;
                    6: level_vec_out = 64'b1011111001111110011010100100011110101110110100001001000100101101;
                    7: level_vec_out = 64'b1011111001111110011010100100011110101110110100001001000100101111;
                    8: level_vec_out = 64'b1011111001111110011010101100011110101110110100001001000100101111;
                    9: level_vec_out = 64'b1011111001111110011010101100011110101110110100001001000100101111;
                    10: level_vec_out = 64'b1011111001111110011010101100011110101110110100001101000100111111;
                    11: level_vec_out = 64'b1011111001111110011010101100011110101110110100001101000100111111;
                    12: level_vec_out = 64'b1011111001111110011010101100011110101110110110001101000100111111;
                    13: level_vec_out = 64'b1011111001111110011010111100011110101110110111001101000100111111;
                    14: level_vec_out = 64'b1011111001111110011010111100111110101111110111001101000100111111;
                    15: level_vec_out = 64'b1011111001111110011010111100111110101111110111001101000101111111;
                    16: level_vec_out = 64'b1011111001111110011011111100111110111111110111001101000101111111;
                    17: level_vec_out = 64'b1011111011111110011011111101111110111111110111001101000101111111;
                    18: level_vec_out = 64'b1011111011111110011011111101111110111111110111011101000101111111;
                    19: level_vec_out = 64'b1011111111111110011011111101111111111111110111011101000101111111;
                    20: level_vec_out = 64'b1011111111111110011011111101111111111111110111011101000101111111;
                    21: level_vec_out = 64'b1011111111111110011011111101111111111111110111111101100101111111;
                    22: level_vec_out = 64'b1011111111111110011111111101111111111111110111111101110101111111;
                    23: level_vec_out = 64'b1011111111111110011111111101111111111111110111111101110101111111;
                    24: level_vec_out = 64'b1011111111111110111111111101111111111111110111111101110101111111;
                    25: level_vec_out = 64'b1011111111111110111111111101111111111111110111111101110101111111;
                    26: level_vec_out = 64'b1011111111111110111111111101111111111111110111111101110101111111;
                    27: level_vec_out = 64'b1011111111111110111111111101111111111111110111111101110101111111;
                    28: level_vec_out = 64'b1011111111111110111111111101111111111111111111111101111111111111;
                    29: level_vec_out = 64'b1011111111111110111111111111111111111111111111111101111111111111;
                    30: level_vec_out = 64'b1011111111111111111111111111111111111111111111111101111111111111;
                    31: level_vec_out = 64'b1011111111111111111111111111111111111111111111111111111111111111;
                endcase
            end
            3: begin
                case (frame_id)
                    0: level_vec_out = 64'b1101010011010000000100111001111001011111100010111101001110111111;
                    1: level_vec_out = 64'b1101010011010000000100111001111001011111100010111101001110111111;
                    2: level_vec_out = 64'b1101010011010000000110111001111001011111100010111101001110111111;
                    3: level_vec_out = 64'b1101010011010000000110111001111001011111100110111101001110111111;
                    4: level_vec_out = 64'b1101010011010000010110111001111001011111100110111101001110111111;
                    5: level_vec_out = 64'b1101010011010000010110111001111001011111100110111101001110111111;
                    6: level_vec_out = 64'b1101010011010100010110111001111001011111100110111101001110111111;
                    7: level_vec_out = 64'b1101010011010100010110111101111001111111100110111101101110111111;
                    8: level_vec_out = 64'b1101010011010100010110111101111001111111100110111101101110111111;
                    9: level_vec_out = 64'b1101110011010100010110111101111001111111100110111101101110111111;
                    10: level_vec_out = 64'b1101110011010100010110111101111001111111100110111101101110111111;
                    11: level_vec_out = 64'b1101110011010100110110111101111001111111100110111111101110111111;
                    12: level_vec_out = 64'b1101110011010100110110111101111001111111100110111111101110111111;
                    13: level_vec_out = 64'b1101110011010100110110111101111001111111100110111111101110111111;
                    14: level_vec_out = 64'b1101110111010100110110111101111001111111100110111111101110111111;
                    15: level_vec_out = 64'b1101110111010100110110111101111001111111100110111111101110111111;
                    16: level_vec_out = 64'b1101110111010100110110111101111001111111100110111111101110111111;
                    17: level_vec_out = 64'b1101110111010100110110111101111001111111100110111111101110111111;
                    18: level_vec_out = 64'b1101110111010100110110111101111001111111100110111111101110111111;
                    19: level_vec_out = 64'b1101110111010100110110111101111001111111110110111111101110111111;
                    20: level_vec_out = 64'b1101111111010100111110111101111001111111110110111111101110111111;
                    21: level_vec_out = 64'b1101111111010100111110111101111001111111110110111111101110111111;
                    22: level_vec_out = 64'b1101111111010100111111111101111001111111110110111111101111111111;
                    23: level_vec_out = 64'b1101111111010100111111111101111001111111110110111111111111111111;
                    24: level_vec_out = 64'b1111111111010100111111111101111101111111110110111111111111111111;
                    25: level_vec_out = 64'b1111111111010110111111111101111101111111111110111111111111111111;
                    26: level_vec_out = 64'b1111111111010110111111111111111111111111111110111111111111111111;
                    27: level_vec_out = 64'b1111111111010111111111111111111111111111111110111111111111111111;
                    28: level_vec_out = 64'b1111111111010111111111111111111111111111111110111111111111111111;
                    29: level_vec_out = 64'b1111111111111111111111111111111111111111111110111111111111111111;
                    30: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    31: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                endcase
            end
            4: begin
                case (frame_id)
                    0: level_vec_out = 64'b1100011001101101000010101110011001011001101100110110111011010001;
                    1: level_vec_out = 64'b1100011001101101000010101110011001011001101100110111111011010001;
                    2: level_vec_out = 64'b1100011001101101000010101110011001011001101100110111111011010001;
                    3: level_vec_out = 64'b1100011001101101000010101110011101011001101100110111111011010001;
                    4: level_vec_out = 64'b1100011001101101000010101110011111011001101100110111111011010001;
                    5: level_vec_out = 64'b1100111001101101000010101110011111011001101100110111111011010001;
                    6: level_vec_out = 64'b1100111001101101000010101110011111011001101100110111111011010001;
                    7: level_vec_out = 64'b1100111001101101000010101110011111011001101100110111111011010101;
                    8: level_vec_out = 64'b1100111001101101001010101110011111011001101100110111111011010101;
                    9: level_vec_out = 64'b1100111111101101001010101110011111011001101110110111111011010101;
                    10: level_vec_out = 64'b1100111111101101001010101110011111011001101110110111111111010101;
                    11: level_vec_out = 64'b1100111111101101001010101110011111011001101110110111111111010101;
                    12: level_vec_out = 64'b1100111111101101001010101110011111011001101110110111111111010101;
                    13: level_vec_out = 64'b1110111111101101001010101110011111011001101110110111111111010101;
                    14: level_vec_out = 64'b1110111111101101001010101110011111011001101110110111111111010101;
                    15: level_vec_out = 64'b1110111111101111011010101110011111011001101110110111111111010101;
                    16: level_vec_out = 64'b1110111111101111011010101110011111011011101110110111111111010101;
                    17: level_vec_out = 64'b1110111111101111011010111110011111011011101110110111111111010101;
                    18: level_vec_out = 64'b1110111111101111011010111110011111011011101110110111111111010111;
                    19: level_vec_out = 64'b1110111111101111011010111110011111011011101110110111111111011111;
                    20: level_vec_out = 64'b1110111111101111011010111110011111111011101110110111111111011111;
                    21: level_vec_out = 64'b1110111111101111011010111110011111111011101110110111111111011111;
                    22: level_vec_out = 64'b1110111111101111011010111111011111111011101111110111111111011111;
                    23: level_vec_out = 64'b1110111111101111011011111111011111111011101111110111111111011111;
                    24: level_vec_out = 64'b1110111111101111011011111111011111111011101111110111111111011111;
                    25: level_vec_out = 64'b1110111111101111011011111111011111111011101111110111111111011111;
                    26: level_vec_out = 64'b1110111111101111011011111111111111111011111111110111111111011111;
                    27: level_vec_out = 64'b1110111111101111011011111111111111111111111111110111111111011111;
                    28: level_vec_out = 64'b1110111111111111011011111111111111111111111111110111111111011111;
                    29: level_vec_out = 64'b1110111111111111011011111111111111111111111111110111111111011111;
                    30: level_vec_out = 64'b1110111111111111111011111111111111111111111111111111111111011111;
                    31: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111011111;
                endcase
            end
            5: begin
                case (frame_id)
                    0: level_vec_out = 64'b0011011111001000100101000000010011011110100001101010100100011100;
                    1: level_vec_out = 64'b0011011111001000100101000000010011011110100101101010100100011100;
                    2: level_vec_out = 64'b0011011111001000100101000000010011011110100101101010110100011100;
                    3: level_vec_out = 64'b0011011111001000100101000000010011011110100101101010110100011100;
                    4: level_vec_out = 64'b0011011111001000100101000000010011011110100101101110110100011100;
                    5: level_vec_out = 64'b0011011111001000100101000000010011011110100101101110110100011100;
                    6: level_vec_out = 64'b0011011111001000100101000000010011011110100101101110110100011100;
                    7: level_vec_out = 64'b0011011111001000100101000000010011111110100101101110110100011100;
                    8: level_vec_out = 64'b0011011111001000100101000000010011111110100101101110110100011100;
                    9: level_vec_out = 64'b0011011111001000100101000000010011111110100101101110110100011100;
                    10: level_vec_out = 64'b0011011111001000100101001000010011111110100101101110110100011100;
                    11: level_vec_out = 64'b0011011111001000100101001000011011111110100101101110111100011100;
                    12: level_vec_out = 64'b0011011111001000101101001100011011111110100101101110111100011100;
                    13: level_vec_out = 64'b0011011111001000101101001100011011111110100101101110111100011100;
                    14: level_vec_out = 64'b0011011111001000101101011100011011111110100101101110111100011100;
                    15: level_vec_out = 64'b0011111111001000101101011100111011111110100101101110111100111100;
                    16: level_vec_out = 64'b0011111111001001101101011100111011111110100101101110111100111100;
                    17: level_vec_out = 64'b0011111111001001101101011110111011111110100101101110111100111101;
                    18: level_vec_out = 64'b0011111111101001101101011110111011111110110101101110111110111101;
                    19: level_vec_out = 64'b0011111111101001101101011110111011111110110101101110111110111101;
                    20: level_vec_out = 64'b0011111111101001111101011110111111111110110101101110111110111101;
                    21: level_vec_out = 64'b0011111111111001111111111110111111111110110101101110111110111101;
                    22: level_vec_out = 64'b0011111111111001111111111110111111111110110101101110111110111111;
                    23: level_vec_out = 64'b0011111111111001111111111110111111111110110101101110111110111111;
                    24: level_vec_out = 64'b0011111111111011111111111110111111111110110101101110111111111111;
                    25: level_vec_out = 64'b0011111111111011111111111110111111111111110111101110111111111111;
                    26: level_vec_out = 64'b0011111111111011111111111111111111111111110111101110111111111111;
                    27: level_vec_out = 64'b1011111111111011111111111111111111111111110111101111111111111111;
                    28: level_vec_out = 64'b1011111111111011111111111111111111111111110111101111111111111111;
                    29: level_vec_out = 64'b1011111111111011111111111111111111111111110111101111111111111111;
                    30: level_vec_out = 64'b1011111111111011111111111111111111111111110111101111111111111111;
                    31: level_vec_out = 64'b1111111111111011111111111111111111111111111111101111111111111111;
                endcase
            end
            6: begin
                case (frame_id)
                    0: level_vec_out = 64'b0101111100101101000111010101111010001111101000001010000011100100;
                    1: level_vec_out = 64'b0101111100101101000111010101111010011111101000001110000011100100;
                    2: level_vec_out = 64'b0101111100101101000111010101111010011111101000001110000011100100;
                    3: level_vec_out = 64'b0101111100101101000111010101111010011111101000001110000011100100;
                    4: level_vec_out = 64'b0111111100101101000111010101111011011111101000001110000011100100;
                    5: level_vec_out = 64'b0111111100101101000111011101111011011111101000001110000011100100;
                    6: level_vec_out = 64'b0111111100101101000111011101111011011111101000001110100111100110;
                    7: level_vec_out = 64'b0111111100101101000111011101111011011111101000001110100111100110;
                    8: level_vec_out = 64'b0111111100101101000111011101111011011111101000001110100111100110;
                    9: level_vec_out = 64'b0111111111101101000111011101111011011111101010001110100111100110;
                    10: level_vec_out = 64'b0111111111101101000111011101111011011111101010001110100111110110;
                    11: level_vec_out = 64'b0111111111101101000111011101111011011111101010001110100111111110;
                    12: level_vec_out = 64'b0111111111101101000111011111111011011111111010001110100111111110;
                    13: level_vec_out = 64'b0111111111101101000111011111111011011111111011001110100111111110;
                    14: level_vec_out = 64'b0111111111101101000111011111111011011111111011001110100111111110;
                    15: level_vec_out = 64'b0111111111101101000111011111111011011111111011001110100111111110;
                    16: level_vec_out = 64'b0111111111101101000111011111111011011111111011001110100111111111;
                    17: level_vec_out = 64'b0111111111101101011111011111111011011111111011001110100111111111;
                    18: level_vec_out = 64'b0111111111101101011111011111111011011111111011001110100111111111;
                    19: level_vec_out = 64'b1111111111101101011111111111111011011111111011001110100111111111;
                    20: level_vec_out = 64'b1111111111101101011111111111111011011111111011001110100111111111;
                    21: level_vec_out = 64'b1111111111101101011111111111111011011111111011001110100111111111;
                    22: level_vec_out = 64'b1111111111101101011111111111111011011111111011001110100111111111;
                    23: level_vec_out = 64'b1111111111101101011111111111111011011111111011001110100111111111;
                    24: level_vec_out = 64'b1111111111101101011111111111111011011111111111001110100111111111;
                    25: level_vec_out = 64'b1111111111101101011111111111111011011111111111001110100111111111;
                    26: level_vec_out = 64'b1111111111101101011111111111111011111111111111001110100111111111;
                    27: level_vec_out = 64'b1111111111101101011111111111111011111111111111111110100111111111;
                    28: level_vec_out = 64'b1111111111111101011111111111111011111111111111111110100111111111;
                    29: level_vec_out = 64'b1111111111111111111111111111111011111111111111111110101111111111;
                    30: level_vec_out = 64'b1111111111111111111111111111111011111111111111111110101111111111;
                    31: level_vec_out = 64'b1111111111111111111111111111111011111111111111111111111111111111;
                endcase
            end
            7: begin
                case (frame_id)
                    0: level_vec_out = 64'b0011011011100110111011100000010101111001111000010010100111010110;
                    1: level_vec_out = 64'b0011011011100110111011100010010101111001111000010010100111010110;
                    2: level_vec_out = 64'b0011011011100110111011100010010101111001111000010010101111010110;
                    3: level_vec_out = 64'b0011011011101110111011100010010101111101111000110010101111010110;
                    4: level_vec_out = 64'b0011011011101110111011100010010101111101111001110010101111010110;
                    5: level_vec_out = 64'b0011011011101110111011100010010101111101111001111010101111010110;
                    6: level_vec_out = 64'b0111011011101111111011100010010101111101111001111010101111010110;
                    7: level_vec_out = 64'b0111111011101111111011100010010101111101111001111010101111010110;
                    8: level_vec_out = 64'b0111111111111111111011100010010101111101111001111010101111010110;
                    9: level_vec_out = 64'b0111111111111111111011100010011101111101111001111010101111010110;
                    10: level_vec_out = 64'b0111111111111111111011100010011101111101111001111010101111010110;
                    11: level_vec_out = 64'b0111111111111111111011110010011101111101111001111010101111010110;
                    12: level_vec_out = 64'b1111111111111111111011110010011101111101111001111010101111010110;
                    13: level_vec_out = 64'b1111111111111111111011110110011101111101111001111010101111010110;
                    14: level_vec_out = 64'b1111111111111111111011110110011101111101111001111010101111010110;
                    15: level_vec_out = 64'b1111111111111111111011110111011101111101111001111010101111010110;
                    16: level_vec_out = 64'b1111111111111111111011110111011101111101111001111110101111010110;
                    17: level_vec_out = 64'b1111111111111111111011110111011101111101111001111110101111010110;
                    18: level_vec_out = 64'b1111111111111111111011110111011101111101111001111110101111010110;
                    19: level_vec_out = 64'b1111111111111111111011110111011101111101111001111110101111010110;
                    20: level_vec_out = 64'b1111111111111111111011110111011101111111111001111110101111010110;
                    21: level_vec_out = 64'b1111111111111111111011110111111101111111111001111110101111010110;
                    22: level_vec_out = 64'b1111111111111111111011110111111101111111111001111110101111010110;
                    23: level_vec_out = 64'b1111111111111111111011110111111111111111111111111110101111110110;
                    24: level_vec_out = 64'b1111111111111111111011110111111111111111111111111110101111110110;
                    25: level_vec_out = 64'b1111111111111111111011110111111111111111111111111110111111110110;
                    26: level_vec_out = 64'b1111111111111111111011110111111111111111111111111110111111111110;
                    27: level_vec_out = 64'b1111111111111111111011110111111111111111111111111110111111111110;
                    28: level_vec_out = 64'b1111111111111111111011111111111111111111111111111110111111111111;
                    29: level_vec_out = 64'b1111111111111111111011111111111111111111111111111111111111111111;
                    30: level_vec_out = 64'b1111111111111111111011111111111111111111111111111111111111111111;
                    31: level_vec_out = 64'b1111111111111111111011111111111111111111111111111111111111111111;
                endcase
            end
        endcase
    end
endmodule