----
 -- @file level_hvec_gen_hdl.hpp
 -- @brief This script generates HDL code for generating high-dimensional LEVEL vectors.
 -- It is a novel method; for more information, please refer to our paper.
 --
 -- @author Saeid Jamili and Marco Angioli
 -- @note Author names are listed in alphabetical order.
 -- @email <saeid.jamili@uniroma1.it>
 -- @email <marco.angioli@uniroma1.it>
 --
 -- @contributors
 --
 -- @date Created: 24th July 2023
 -- @date Last Updated: 23th August 2023
 --
 -- @version 1.0.0
 --
 -- @institute Sapienza University of Rome
 -- @cite https://doi.org/10.xxxx/yyyyy
 --
 -- @section DEPENDENCIES
 -- - Dependency1: Description or version details.
 -- - Dependency2: Description or version details.
 --
 -- @section LICENSE
 -- This file is part of the Aeneas HyperCompute Platform.
 --
 -- Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 --
 -- @section CHANGELOG
 -- @version 1.0.0-dev - 23th August 2023
 -- - Initial release
 --
 -- @todo
 -- - Complete level vector generator function
 -- - Add training
 --
 -- @see
 -- -
 -- -
 -- -
 --
 --

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity level_vec_gen is
    Port ( level_vec_out : out  STD_LOGIC_VECTOR (63 downto 0);
           frame_index : in  STD_LOGIC_VECTOR (2 downto 0);
           frame_id : in  STD_LOGIC_VECTOR (4 downto 0));
end level_vec_gen;

architecture Behavioral of level_vec_gen is
begin
    process (frame_index, frame_id)
    begin
        -- Update this function to match your requirements
        case frame_index is
            when "000" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1100100101000110000111011100101011100001111000000111010110000110";
                    when "00001" => level_vec_out <= "1100100101000110010111011100101011100001111000000111010110001110";
                    when "00010" => level_vec_out <= "1100100101000110011111011100101011100001111010000111011110001110";
                    when "00011" => level_vec_out <= "1100100101000110011111011100101011100001111011000111011110001110";
                    when "00100" => level_vec_out <= "1100100101000110011111011100101011100001111011000111011110001110";
                    when "00101" => level_vec_out <= "1110100101000110011111011100101011100001111011000111011110001110";
                    when "00110" => level_vec_out <= "1110100101000110011111011100101011100001111011000111011110001110";
                    when "00111" => level_vec_out <= "1110100101000110011111111100101011100001111011000111011110001110";
                    when "01000" => level_vec_out <= "1110100101000110011111111100101111100001111011000111011110001110";
                    when "01001" => level_vec_out <= "1110100101000110011111111100101111100001111011000111011110001110";
                    when "01010" => level_vec_out <= "1110100101000110011111111100101111110001111011000111011110001110";
                    when "01011" => level_vec_out <= "1110100101000110011111111100101111110001111011000111011110001110";
                    when "01100" => level_vec_out <= "1110100101000110011111111100101111110001111011010111011110011110";
                    when "01101" => level_vec_out <= "1110100111000110111111111100101111111001111011010111011110011110";
                    when "01110" => level_vec_out <= "1110101111000110111111111100101111111001111011110111011110011110";
                    when "01111" => level_vec_out <= "1110101111000110111111111100101111111001111011111111011110111110";
                    when "10000" => level_vec_out <= "1110101111010110111111111100101111111001111011111111011110111110";
                    when "10001" => level_vec_out <= "1110101111110110111111111100101111111001111011111111011110111110";
                    when "10010" => level_vec_out <= "1110101111110110111111111100101111111001111011111111011110111110";
                    when "10011" => level_vec_out <= "1110101111110110111111111100101111111001111011111111011110111110";
                    when "10100" => level_vec_out <= "1110101111110110111111111100101111111011111011111111011110111110";
                    when "10101" => level_vec_out <= "1110101111110110111111111100101111111011111011111111011111111111";
                    when "10110" => level_vec_out <= "1110101111110110111111111100101111111011111111111111011111111111";
                    when "10111" => level_vec_out <= "1110111111110110111111111100101111111011111111111111011111111111";
                    when "11000" => level_vec_out <= "1110111111110110111111111110111111111011111111111111011111111111";
                    when "11001" => level_vec_out <= "1110111111110110111111111110111111111011111111111111011111111111";
                    when "11010" => level_vec_out <= "1110111111110110111111111110111111111011111111111111011111111111";
                    when "11011" => level_vec_out <= "1110111111110110111111111111111111111011111111111111011111111111";
                    when "11100" => level_vec_out <= "1110111111110110111111111111111111111011111111111111011111111111";
                    when "11101" => level_vec_out <= "1110111111110110111111111111111111111011111111111111011111111111";
                    when "11110" => level_vec_out <= "1111111111111110111111111111111111111011111111111111011111111111";
                    when "11111" => level_vec_out <= "1111111111111110111111111111111111111011111111111111011111111111";
                when others => null;
                end case;
            when "001" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0011011100100010111101010110001011001111100110110101000111010010";
                    when "00001" => level_vec_out <= "0011011100100010111101010110001011001111100110110101000111010010";
                    when "00010" => level_vec_out <= "0011011100100010111101010110001011001111100110110101000111010010";
                    when "00011" => level_vec_out <= "0011011100100011111101010111001011001111101110110101001111010010";
                    when "00100" => level_vec_out <= "0011011100100011111101010111001011001111101110110101001111010010";
                    when "00101" => level_vec_out <= "0011011100100011111101010111001011001111101110110101001111010010";
                    when "00110" => level_vec_out <= "0011011100100011111101010111001011001111101110110101101111010010";
                    when "00111" => level_vec_out <= "0011011100100011111101010111001011001111101110110101101111010010";
                    when "01000" => level_vec_out <= "0011011100100011111101110111001011001111101111110101101111010110";
                    when "01001" => level_vec_out <= "0011011100100011111101110111001011001111101111110101101111010110";
                    when "01010" => level_vec_out <= "0011011100100011111101110111011011001111101111110101101111010110";
                    when "01011" => level_vec_out <= "0011011100100011111101111111011111001111101111110101101111010110";
                    when "01100" => level_vec_out <= "0011111100100011111101111111011111001111101111111101101111010110";
                    when "01101" => level_vec_out <= "0011111100100011111101111111011111001111101111111101101111010110";
                    when "01110" => level_vec_out <= "0011111100100011111101111111011111001111101111111101101111110110";
                    when "01111" => level_vec_out <= "0011111100110011111101111111011111011111101111111101101111110110";
                    when "10000" => level_vec_out <= "0011111100110011111101111111111111011111101111111101101111110110";
                    when "10001" => level_vec_out <= "0011111100110011111101111111111111011111101111111101101111110110";
                    when "10010" => level_vec_out <= "0011111100110011111101111111111111011111101111111101101111110110";
                    when "10011" => level_vec_out <= "0011111110110011111101111111111111011111101111111101101111110110";
                    when "10100" => level_vec_out <= "0011111110110011111101111111111111011111101111111101101111110110";
                    when "10101" => level_vec_out <= "0011111110110011111111111111111111011111101111111101101111110111";
                    when "10110" => level_vec_out <= "0011111110110011111111111111111111011111101111111111101111110111";
                    when "10111" => level_vec_out <= "0011111110111011111111111111111111011111101111111111101111110111";
                    when "11000" => level_vec_out <= "0011111110111011111111111111111111011111101111111111101111110111";
                    when "11001" => level_vec_out <= "0111111110111011111111111111111111011111111111111111101111110111";
                    when "11010" => level_vec_out <= "1111111111111011111111111111111111011111111111111111101111111111";
                    when "11011" => level_vec_out <= "1111111111111011111111111111111111011111111111111111111111111111";
                    when "11100" => level_vec_out <= "1111111111111011111111111111111111011111111111111111111111111111";
                    when "11101" => level_vec_out <= "1111111111111011111111111111111111111111111111111111111111111111";
                    when "11110" => level_vec_out <= "1111111111111011111111111111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "010" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1100110111001010101100110100000001111010001011110101011110000110";
                    when "00001" => level_vec_out <= "1100110111001010101110110100000001111010001011110101011110000110";
                    when "00010" => level_vec_out <= "1100110111001010101110110100000001111010001011110101011110000110";
                    when "00011" => level_vec_out <= "1100110111001010101110110100000011111010001011110101011110000110";
                    when "00100" => level_vec_out <= "1100110111011010101110110110000011111010001011110101011110000110";
                    when "00101" => level_vec_out <= "1100110111011010101110110110000011111110001011110101011110000110";
                    when "00110" => level_vec_out <= "1100110111011010111110110110000011111110001011110101011110010110";
                    when "00111" => level_vec_out <= "1100111111011010111110110110000011111110001011110101011110010110";
                    when "01000" => level_vec_out <= "1100111111011010111111110110000011111110001011110101011110010110";
                    when "01001" => level_vec_out <= "1100111111011010111111110110000011111110101011110101011110010110";
                    when "01010" => level_vec_out <= "1100111111011010111111110110000011111110101011110101011110010110";
                    when "01011" => level_vec_out <= "1100111111111010111111110110000011111110101011110101111110010110";
                    when "01100" => level_vec_out <= "1100111111111010111111110110000011111110101011110101111110010110";
                    when "01101" => level_vec_out <= "1100111111111010111111110110010011111111101111110101111110010110";
                    when "01110" => level_vec_out <= "1110111111111010111111110110010011111111101111110101111110010110";
                    when "01111" => level_vec_out <= "1110111111111010111111110110010011111111101111110101111110010110";
                    when "10000" => level_vec_out <= "1110111111111010111111111110010011111111111111110101111110010110";
                    when "10001" => level_vec_out <= "1111111111111011111111111110010011111111111111110101111110011110";
                    when "10010" => level_vec_out <= "1111111111111011111111111110010011111111111111110101111110011110";
                    when "10011" => level_vec_out <= "1111111111111011111111111111010011111111111111110101111110011110";
                    when "10100" => level_vec_out <= "1111111111111011111111111111110011111111111111110101111110011110";
                    when "10101" => level_vec_out <= "1111111111111011111111111111110011111111111111110101111110011110";
                    when "10110" => level_vec_out <= "1111111111111011111111111111110011111111111111110101111110011110";
                    when "10111" => level_vec_out <= "1111111111111011111111111111110111111111111111110101111111011110";
                    when "11000" => level_vec_out <= "1111111111111011111111111111110111111111111111110101111111011110";
                    when "11001" => level_vec_out <= "1111111111111011111111111111110111111111111111110111111111011110";
                    when "11010" => level_vec_out <= "1111111111111011111111111111110111111111111111110111111111011111";
                    when "11011" => level_vec_out <= "1111111111111011111111111111110111111111111111110111111111111111";
                    when "11100" => level_vec_out <= "1111111111111011111111111111110111111111111111111111111111111111";
                    when "11101" => level_vec_out <= "1111111111111011111111111111110111111111111111111111111111111111";
                    when "11110" => level_vec_out <= "1111111111111011111111111111110111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111011111111111111110111111111111111111111111111111111";
                when others => null;
                end case;
            when "011" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0010001000100101011111100010100010001010101001110100111010110100";
                    when "00001" => level_vec_out <= "0011001000100101111111100010100010001010101001110100111010110100";
                    when "00010" => level_vec_out <= "0011001000100101111111100010100010001010101001110100111010110100";
                    when "00011" => level_vec_out <= "0011001000100101111111100010100010001010101001110100111010110100";
                    when "00100" => level_vec_out <= "0011001000100101111111100010100110001010101011110100111010110100";
                    when "00101" => level_vec_out <= "0011001000100101111111100010100110001010101011110100111010110100";
                    when "00110" => level_vec_out <= "0011011000100101111111100010100110001010101011110100111010110100";
                    when "00111" => level_vec_out <= "0011011000100111111111100010100110001010101011110100111010110100";
                    when "01000" => level_vec_out <= "0011011001101111111111100010100110001010101011110100111010110100";
                    when "01001" => level_vec_out <= "0011011001101111111111100010100110001010101011111100111010110100";
                    when "01010" => level_vec_out <= "0011011001101111111111100010100110001010101011111100111110110100";
                    when "01011" => level_vec_out <= "0011011001101111111111100010100110001010101011111100111110110100";
                    when "01100" => level_vec_out <= "0011011001101111111111100010100110001010101011111100111110110100";
                    when "01101" => level_vec_out <= "0011011001101111111111100010100110001010101011111100111110110100";
                    when "01110" => level_vec_out <= "0011011001101111111111100010100110001010111011111100111110110100";
                    when "01111" => level_vec_out <= "0011011001101111111111100010100110001010111011111100111110110100";
                    when "10000" => level_vec_out <= "1011011001101111111111100110100110001010111011111100111110110100";
                    when "10001" => level_vec_out <= "1011011001101111111111100110100110001010111011111100111110110100";
                    when "10010" => level_vec_out <= "1011011001101111111111110110110110001010111011111100111110111100";
                    when "10011" => level_vec_out <= "1011011001101111111111110111110110001010111011111100111110111100";
                    when "10100" => level_vec_out <= "1011011001101111111111110111110110101010111011111100111111111110";
                    when "10101" => level_vec_out <= "1011011101101111111111110111110110101010111011111100111111111110";
                    when "10110" => level_vec_out <= "1011111101101111111111110111110110101010111011111100111111111111";
                    when "10111" => level_vec_out <= "1011111101101111111111110111110110101010111011111100111111111111";
                    when "11000" => level_vec_out <= "1011111111101111111111111111110110101010111011111100111111111111";
                    when "11001" => level_vec_out <= "1011111111101111111111111111110110101010111111111100111111111111";
                    when "11010" => level_vec_out <= "1111111111101111111111111111110110101010111111111100111111111111";
                    when "11011" => level_vec_out <= "1111111111101111111111111111110110111110111111111100111111111111";
                    when "11100" => level_vec_out <= "1111111111101111111111111111110110111110111111111100111111111111";
                    when "11101" => level_vec_out <= "1111111111101111111111111111110110111110111111111101111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111110111111110111111111101111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "100" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0011010000100011101101010010010100111100111000101101110100011010";
                    when "00001" => level_vec_out <= "0011010000100011101101010010011100111100111000101101110100011010";
                    when "00010" => level_vec_out <= "1011010000100011101101010010011100111100111000111101110100011010";
                    when "00011" => level_vec_out <= "1011010000100011101101010010011100111100111000111101110100011010";
                    when "00100" => level_vec_out <= "1011010000100011101101010010011100111100111000111101110100011011";
                    when "00101" => level_vec_out <= "1011010001100011101101010010011110111100111000111101110100011011";
                    when "00110" => level_vec_out <= "1011010001100011101101010010011110111100111000111101110100011011";
                    when "00111" => level_vec_out <= "1111010001110011101101010010011110111100111000111101110100011011";
                    when "01000" => level_vec_out <= "1111010001110011101101010010011110111100111000111101110100011011";
                    when "01001" => level_vec_out <= "1111010011110011101101010010011110111100111001111101110100011011";
                    when "01010" => level_vec_out <= "1111010011110011101101010010011110111100111001111101110100011011";
                    when "01011" => level_vec_out <= "1111010011110011101101010010011110111100111001111101110100011011";
                    when "01100" => level_vec_out <= "1111010011110011101101011010011111111100111001111101110100011011";
                    when "01101" => level_vec_out <= "1111010011111011101101011010011111111100111001111101110100011011";
                    when "01110" => level_vec_out <= "1111010011111011101101011010011111111100111001111101110100011011";
                    when "01111" => level_vec_out <= "1111011011111011101101011011011111111100111001111101110101011011";
                    when "10000" => level_vec_out <= "1111011011111011101101011011011111111100111001111101110101111011";
                    when "10001" => level_vec_out <= "1111111011111011101101011011011111111100111001111101110101111011";
                    when "10010" => level_vec_out <= "1111111011111011101101011011011111111100111001111101110101111011";
                    when "10011" => level_vec_out <= "1111111011111011101101011011011111111110111101111101110101111011";
                    when "10100" => level_vec_out <= "1111111011111011101101011011011111111110111101111101110101111011";
                    when "10101" => level_vec_out <= "1111111011111011101101011011011111111110111101111101110101111011";
                    when "10110" => level_vec_out <= "1111111111111011101101011011011111111110111101111101110111111011";
                    when "10111" => level_vec_out <= "1111111111111011101101011011011111111110111101111111110111111111";
                    when "11000" => level_vec_out <= "1111111111111011101101011111011111111110111101111111110111111111";
                    when "11001" => level_vec_out <= "1111111111111011101101011111011111111111111111111111110111111111";
                    when "11010" => level_vec_out <= "1111111111111011111111011111011111111111111111111111110111111111";
                    when "11011" => level_vec_out <= "1111111111111011111111011111011111111111111111111111110111111111";
                    when "11100" => level_vec_out <= "1111111111111011111111011111111111111111111111111111110111111111";
                    when "11101" => level_vec_out <= "1111111111111111111111011111111111111111111111111111110111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "101" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0011101111100001110001010100000100001110100001011011101001101011";
                    when "00001" => level_vec_out <= "0011101111100001110001011100000100001110100001011011101001101011";
                    when "00010" => level_vec_out <= "0011101111100001110001011100000100001110100001111011101001101011";
                    when "00011" => level_vec_out <= "0011111111100001110001011100000100001110100001111011101001101011";
                    when "00100" => level_vec_out <= "0011111111100001110001011100000100001110100001111011101001101011";
                    when "00101" => level_vec_out <= "0011111111100001110001011100000100001110100001111011101001101011";
                    when "00110" => level_vec_out <= "0011111111100101110001011100001100001111100001111011101001101011";
                    when "00111" => level_vec_out <= "0011111111100101110001011100001100011111100001111011101001101011";
                    when "01000" => level_vec_out <= "0011111111100101110001011100001100011111100001111011101001101011";
                    when "01001" => level_vec_out <= "0011111111100101110001011100101100011111100001111011101001101011";
                    when "01010" => level_vec_out <= "0011111111100101110001011100101101011111100001111111111001101011";
                    when "01011" => level_vec_out <= "0011111111100101110001011100101111011111100001111111111001101011";
                    when "01100" => level_vec_out <= "0011111111100101110001011100101111011111100001111111111001101011";
                    when "01101" => level_vec_out <= "0011111111100101110001011100101111011111100001111111111001101011";
                    when "01110" => level_vec_out <= "0011111111100101110001011100111111011111100001111111111001101011";
                    when "01111" => level_vec_out <= "0011111111100101110001011100111111011111100001111111111001101011";
                    when "10000" => level_vec_out <= "0011111111100101110001011100111111011111100001111111111001101011";
                    when "10001" => level_vec_out <= "0011111111100101110001111100111111011111100001111111111001101011";
                    when "10010" => level_vec_out <= "0111111111101101110101111100111111011111100001111111111001101011";
                    when "10011" => level_vec_out <= "0111111111101101110101111100111111011111100001111111111001101111";
                    when "10100" => level_vec_out <= "0111111111101101110101111110111111011111110001111111111001101111";
                    when "10101" => level_vec_out <= "0111111111101101111111111110111111011111110001111111111001101111";
                    when "10110" => level_vec_out <= "1111111111101101111111111110111111011111110001111111111001101111";
                    when "10111" => level_vec_out <= "1111111111101101111111111111111111011111110001111111111001101111";
                    when "11000" => level_vec_out <= "1111111111101101111111111111111111011111110001111111111001101111";
                    when "11001" => level_vec_out <= "1111111111101101111111111111111111011111110001111111111001101111";
                    when "11010" => level_vec_out <= "1111111111101101111111111111111111011111110001111111111001101111";
                    when "11011" => level_vec_out <= "1111111111101101111111111111111111111111110001111111111001101111";
                    when "11100" => level_vec_out <= "1111111111111101111111111111111111111111110101111111111111101111";
                    when "11101" => level_vec_out <= "1111111111111101111111111111111111111111111111111111111111101111";
                    when "11110" => level_vec_out <= "1111111111111101111111111111111111111111111111111111111111101111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111101111";
                when others => null;
                end case;
            when "110" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1100101000110110111101100010000110110110001001011001011111100111";
                    when "00001" => level_vec_out <= "1100101000110110111101100010000110110110001001011001011111100111";
                    when "00010" => level_vec_out <= "1100101000111110111101100010000110110110001001011001011111100111";
                    when "00011" => level_vec_out <= "1100101000111110111101100010000110110110001001011001011111100111";
                    when "00100" => level_vec_out <= "1100101000111110111101110010000110110110001001011011011111100111";
                    when "00101" => level_vec_out <= "1100101000111110111101110110000110110110001001011011011111100111";
                    when "00110" => level_vec_out <= "1100101000111111111101110110000110110110001001011011011111100111";
                    when "00111" => level_vec_out <= "1100101000111111111101110110000110110110011001011011011111100111";
                    when "01000" => level_vec_out <= "1100101000111111111101110110000110110110011001011011011111100111";
                    when "01001" => level_vec_out <= "1100101010111111111101110110000110110110011001011011011111101111";
                    when "01010" => level_vec_out <= "1100101010111111111101110111000110110110011001011011011111101111";
                    when "01011" => level_vec_out <= "1100101010111111111101110111000111110110011001011011011111101111";
                    when "01100" => level_vec_out <= "1100101010111111111101111111000111110110011001011011011111101111";
                    when "01101" => level_vec_out <= "1100101010111111111101111111000111111110011001011011011111101111";
                    when "01110" => level_vec_out <= "1100101010111111111101111111000111111110011001111011011111101111";
                    when "01111" => level_vec_out <= "1100101010111111111101111111000111111110011001111011011111101111";
                    when "10000" => level_vec_out <= "1100101010111111111101111111000111111110011001111011011111101111";
                    when "10001" => level_vec_out <= "1100101010111111111101111111000111111110011001111011111111101111";
                    when "10010" => level_vec_out <= "1100101110111111111101111111000111111110011101111011111111101111";
                    when "10011" => level_vec_out <= "1100101110111111111101111111001111111110011101111011111111101111";
                    when "10100" => level_vec_out <= "1100101110111111111101111111011111111110011101111011111111101111";
                    when "10101" => level_vec_out <= "1100101110111111111101111111011111111110011101111011111111101111";
                    when "10110" => level_vec_out <= "1100101111111111111101111111011111111110011101111011111111101111";
                    when "10111" => level_vec_out <= "1100101111111111111101111111011111111110011101111011111111101111";
                    when "11000" => level_vec_out <= "1100111111111111111101111111111111111111011101111011111111101111";
                    when "11001" => level_vec_out <= "1100111111111111111101111111111111111111011101111011111111101111";
                    when "11010" => level_vec_out <= "1100111111111111111101111111111111111111011101111011111111101111";
                    when "11011" => level_vec_out <= "1100111111111111111101111111111111111111011101111011111111101111";
                    when "11100" => level_vec_out <= "1100111111111111111101111111111111111111011101111111111111101111";
                    when "11101" => level_vec_out <= "1110111111111111111101111111111111111111111101111111111111111111";
                    when "11110" => level_vec_out <= "1110111111111111111111111111111111111111111101111111111111111111";
                    when "11111" => level_vec_out <= "1110111111111111111111111111111111111111111101111111111111111111";
                when others => null;
                end case;
            when "111" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0111000110011011100100011111011111010110100110010110000110000001";
                    when "00001" => level_vec_out <= "0111000110011011100110011111011111010110100110010110000110000001";
                    when "00010" => level_vec_out <= "0111000110011011100110011111011111010111100110010110000110000001";
                    when "00011" => level_vec_out <= "0111000110011011100110011111111111010111100110010110000110000001";
                    when "00100" => level_vec_out <= "0111000110011011100110011111111111010111100110010110000110000011";
                    when "00101" => level_vec_out <= "0111100110111011100111011111111111010111100110010110000110000011";
                    when "00110" => level_vec_out <= "0111100110111011100111011111111111010111100110010110000110000011";
                    when "00111" => level_vec_out <= "0111100110111011100111111111111111010111100110010110000110000011";
                    when "01000" => level_vec_out <= "0111100110111011100111111111111111011111100110010110000110000011";
                    when "01001" => level_vec_out <= "0111100110111011100111111111111111011111100110010110000110000111";
                    when "01010" => level_vec_out <= "0111100110111011100111111111111111111111100110010110000110000111";
                    when "01011" => level_vec_out <= "0111110110111011100111111111111111111111110110010110000110000111";
                    when "01100" => level_vec_out <= "0111111110111011100111111111111111111111110110010110000110000111";
                    when "01101" => level_vec_out <= "0111111110111011100111111111111111111111110110010110000110000111";
                    when "01110" => level_vec_out <= "0111111110111011100111111111111111111111110110110110000110000111";
                    when "01111" => level_vec_out <= "0111111110111011100111111111111111111111110110110110010110000111";
                    when "10000" => level_vec_out <= "1111111110111011100111111111111111111111110110110110010110000111";
                    when "10001" => level_vec_out <= "1111111110111011101111111111111111111111110110110110010110000111";
                    when "10010" => level_vec_out <= "1111111110111011101111111111111111111111110110110110010110000111";
                    when "10011" => level_vec_out <= "1111111110111011111111111111111111111111110110110110010110000111";
                    when "10100" => level_vec_out <= "1111111110111011111111111111111111111111110110110110010110000111";
                    when "10101" => level_vec_out <= "1111111110111011111111111111111111111111110110110110110110000111";
                    when "10110" => level_vec_out <= "1111111110111011111111111111111111111111110110110110110110000111";
                    when "10111" => level_vec_out <= "1111111110111011111111111111111111111111110110110110110111000111";
                    when "11000" => level_vec_out <= "1111111110111011111111111111111111111111110110110110110111000111";
                    when "11001" => level_vec_out <= "1111111111111011111111111111111111111111110110111110110111000111";
                    when "11010" => level_vec_out <= "1111111111111011111111111111111111111111110110111111110111000111";
                    when "11011" => level_vec_out <= "1111111111111011111111111111111111111111110110111111110111011111";
                    when "11100" => level_vec_out <= "1111111111111011111111111111111111111111110110111111111111011111";
                    when "11101" => level_vec_out <= "1111111111111011111111111111111111111111110110111111111111011111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111110110111111111111011111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when others => null;
        end case;
    end process;
end Behavioral;