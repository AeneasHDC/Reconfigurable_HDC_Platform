/**
 * @file level_hvec_gen_hdl.hpp
 * @brief This script generates HDL code for generating high-dimensional LEVEL vectors.
 * It is a novel method; for more information, please refer to our paper.
 *
 * @author Saeid Jamili and Marco Angioli
 * @note Author names are listed in alphabetical order.
 * @email <saeid.jamili@uniroma1.it>
 * @email <marco.angioli@uniroma1.it>
 *
 * @contributors
 *
 * @date Created: 24th July 2023
 * @date Last Updated: 23th August 2023
 *
 * @version 1.0.0
 *
 * @institute Sapienza University of Rome
 * @cite https://doi.org/10.xxxx/yyyyy
 *
 * @section DEPENDENCIES
 * - Dependency1: Description or version details.
 * - Dependency2: Description or version details.
 *
 * @section LICENSE
 * This file is part of the Aeneas HyperCompute Platform.
 *
 * Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 *
 * @section CHANGELOG
 * @version 1.0.0-dev - 23th August 2023
 * - Initial release
 *
 * @todo
 * - Complete level vector generator function
 * - Add training
 *
 * @see
 * -
 * -
 * -
 *
 */

module level_hvec_gen #(parameter int DI_PARALLEL_W_BITS = 64) (
  input logic [2:0] frame_index,
  input logic [4:0] frame_id,
  output logic [DI_PARALLEL_W_BITS-1:0] level_vec_out
);
  always_comb begin
    case (frame_index)
      0:
        case (frame_id)
          0:
            level_vec_out = 64'b0100011100111011010011101100000101011100000110101000111000010000;
          1:
            level_vec_out = 64'b0100011100111011010011101100100101011100001110101000111000010000;
          2:
            level_vec_out = 64'b0100011100111011010011101100100101011100001110111000111000010000;
          3:
            level_vec_out = 64'b0100011100111011010011101100100101011100001110111000111000010000;
          4:
            level_vec_out = 64'b0101011100111011010011101100100101011100001110111000111000010000;
          5:
            level_vec_out = 64'b0101011100111011010111101100100101011100001110111000111000010000;
          6:
            level_vec_out = 64'b0101011100111111010111101100100101011100001110111000111001010001;
          7:
            level_vec_out = 64'b0101011100111111010111101100100101011100001110111000111001010001;
          8:
            level_vec_out = 64'b0101011100111111010111101100100101011100001110111000111101110001;
          9:
            level_vec_out = 64'b0101011100111111010111101100100101111100011110111000111101110001;
          10:
            level_vec_out = 64'b0101011100111111010111101100100101111100011110111000111101110101;
          11:
            level_vec_out = 64'b0101011100111111010111101100100101111100011110111001111101110101;
          12:
            level_vec_out = 64'b0111011100111111010111101110100101111100011110111001111101110101;
          13:
            level_vec_out = 64'b0111011100111111010111101110100101111100011110111001111101110101;
          14:
            level_vec_out = 64'b0111011100111111010111101110100101111110011110111001111101110101;
          15:
            level_vec_out = 64'b0111011100111111010111101110100101111110011110111001111101110101;
          16:
            level_vec_out = 64'b0111011100111111010111101110100101111110011110111001111101110101;
          17:
            level_vec_out = 64'b0111011110111111010111101111100101111111011110111001111101110101;
          18:
            level_vec_out = 64'b1111011110111111010111101111100101111111011111111001111101110101;
          19:
            level_vec_out = 64'b1111011110111111010111101111100101111111011111111001111101110101;
          20:
            level_vec_out = 64'b1111011110111111010111101111100101111111011111111001111101110101;
          21:
            level_vec_out = 64'b1111011110111111010111101111100101111111011111111001111101110101;
          22:
            level_vec_out = 64'b1111111110111111010111101111100101111111011111111001111101110101;
          23:
            level_vec_out = 64'b1111111110111111010111101111100101111111011111111001111101110101;
          24:
            level_vec_out = 64'b1111111110111111010111101111100101111111011111111001111101110101;
          25:
            level_vec_out = 64'b1111111110111111010111101111100101111111011111111001111101111111;
          26:
            level_vec_out = 64'b1111111110111111111111101111100101111111011111111001111101111111;
          27:
            level_vec_out = 64'b1111111110111111111111101111100101111111011111111001111101111111;
          28:
            level_vec_out = 64'b1111111111111111111111101111100101111111111111111101111101111111;
          29:
            level_vec_out = 64'b1111111111111111111111101111110101111111111111111101111111111111;
          30:
            level_vec_out = 64'b1111111111111111111111101111111111111111111111111101111111111111;
          31:
            level_vec_out = 64'b1111111111111111111111101111111111111111111111111111111111111111;
        endcase
      1:
        case (frame_id)
          0:
            level_vec_out = 64'b1110011110001101101111110101101001101111111011101000110010110010;
          1:
            level_vec_out = 64'b1110011110001101101111111101101101101111111011101000110010110010;
          2:
            level_vec_out = 64'b1110011110101101101111111101101101101111111011101000110010110010;
          3:
            level_vec_out = 64'b1110011110101101101111111101101111101111111011101000110010110010;
          4:
            level_vec_out = 64'b1110011110101101101111111101101111101111111011101000110010110110;
          5:
            level_vec_out = 64'b1110011110101101101111111101101111101111111011101000110010110110;
          6:
            level_vec_out = 64'b1110011110101101101111111101101111101111111011101000110010110110;
          7:
            level_vec_out = 64'b1110011110101101101111111101101111101111111011101001110010110110;
          8:
            level_vec_out = 64'b1110011110101101101111111101101111101111111011101001110010110110;
          9:
            level_vec_out = 64'b1110011110101101101111111101101111101111111011101001110010110110;
          10:
            level_vec_out = 64'b1110011110101101101111111101101111101111111011101001110010110110;
          11:
            level_vec_out = 64'b1110011110101101101111111101101111101111111011101001110010110110;
          12:
            level_vec_out = 64'b1110011110101101101111111101101111101111111011101001110011110110;
          13:
            level_vec_out = 64'b1110111110101101101111111101101111101111111011101001110011110110;
          14:
            level_vec_out = 64'b1110111110101101101111111101101111101111111011111001110011110110;
          15:
            level_vec_out = 64'b1110111110101101101111111101101111101111111011111001110011110110;
          16:
            level_vec_out = 64'b1110111110101101111111111101101111101111111011111001110011110110;
          17:
            level_vec_out = 64'b1110111110101101111111111101101111101111111011111001110011110111;
          18:
            level_vec_out = 64'b1110111110101101111111111101101111101111111011111001110011110111;
          19:
            level_vec_out = 64'b1110111110101101111111111101101111101111111011111001110011110111;
          20:
            level_vec_out = 64'b1110111110101101111111111101101111101111111011111001110011110111;
          21:
            level_vec_out = 64'b1110111110101101111111111101101111101111111011111001110111110111;
          22:
            level_vec_out = 64'b1110111110101101111111111101101111101111111011111001110111111111;
          23:
            level_vec_out = 64'b1110111110101111111111111111101111101111111011111001110111111111;
          24:
            level_vec_out = 64'b1110111110101111111111111111101111101111111011111001110111111111;
          25:
            level_vec_out = 64'b1110111110101111111111111111101111111111111011111001110111111111;
          26:
            level_vec_out = 64'b1110111110101111111111111111101111111111111011111001110111111111;
          27:
            level_vec_out = 64'b1110111110101111111111111111101111111111111111111011110111111111;
          28:
            level_vec_out = 64'b1110111110101111111111111111101111111111111111111011110111111111;
          29:
            level_vec_out = 64'b1110111110101111111111111111101111111111111111111011110111111111;
          30:
            level_vec_out = 64'b1111111110101111111111111111101111111111111111111011110111111111;
          31:
            level_vec_out = 64'b1111111110101111111111111111111111111111111111111111110111111111;
        endcase
      2:
        case (frame_id)
          0:
            level_vec_out = 64'b1100110010101000100100101000110011001011011011000100001111101001;
          1:
            level_vec_out = 64'b1100110010101000100100101000110011001011011011000100001111101001;
          2:
            level_vec_out = 64'b1100110010101000100101111001110011001011011011000100001111101001;
          3:
            level_vec_out = 64'b1100110010101000100101111001110011001011011011000100001111101001;
          4:
            level_vec_out = 64'b1100110010101000100101111001110011011011011011000100001111101001;
          5:
            level_vec_out = 64'b1100110010101000100101111001110011011011011011000100001111101101;
          6:
            level_vec_out = 64'b1100110010101000100101111001110011011011011011000100001111101101;
          7:
            level_vec_out = 64'b1100110010101001100101111001110011011011011011000100001111101101;
          8:
            level_vec_out = 64'b1100110010101001100101111001110011011011011011000100011111101101;
          9:
            level_vec_out = 64'b1100110010101001100101111001110011011011011011000100011111101101;
          10:
            level_vec_out = 64'b1100110010101011100101111001111011011011111011000100011111101101;
          11:
            level_vec_out = 64'b1100110010101011100101111001111011011011111011000110011111101101;
          12:
            level_vec_out = 64'b1100110010101011100101111001111011011011111111000111011111101101;
          13:
            level_vec_out = 64'b1100110010101011100101111001111011011011111111000111011111101101;
          14:
            level_vec_out = 64'b1100110010101011100101111001111011011011111111000111011111101101;
          15:
            level_vec_out = 64'b1110110010101011100101111001111011011011111111000111011111101101;
          16:
            level_vec_out = 64'b1110110010101011100101111101111011011011111111001111011111101101;
          17:
            level_vec_out = 64'b1110110010101011100101111101111011011011111111001111011111101101;
          18:
            level_vec_out = 64'b1110110010101011101101111101111011011011111111011111011111101101;
          19:
            level_vec_out = 64'b1110110011111011101101111111111011011011111111011111011111101101;
          20:
            level_vec_out = 64'b1110111011111011101101111111111011011011111111011111011111101101;
          21:
            level_vec_out = 64'b1110111011111011101111111111111011011011111111011111011111101101;
          22:
            level_vec_out = 64'b1110111011111011101111111111111011011011111111011111011111101101;
          23:
            level_vec_out = 64'b1110111011111011101111111111111011111011111111011111011111101101;
          24:
            level_vec_out = 64'b1110111111111011101111111111111011111011111111011111011111101101;
          25:
            level_vec_out = 64'b1111111111111011101111111111111011111011111111011111011111101101;
          26:
            level_vec_out = 64'b1111111111111111101111111111111011111011111111011111011111101111;
          27:
            level_vec_out = 64'b1111111111111111101111111111111011111011111111011111011111111111;
          28:
            level_vec_out = 64'b1111111111111111111111111111111011111011111111011111011111111111;
          29:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111011111011111111111;
          30:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111011111011111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111011111111111;
        endcase
      3:
        case (frame_id)
          0:
            level_vec_out = 64'b0001011001110101101011101010001011101101100111011000100100100011;
          1:
            level_vec_out = 64'b0001111001110101101011101010001011101101100111011000100100100011;
          2:
            level_vec_out = 64'b0001111001110101101011101010001011101101100111011000100100100011;
          3:
            level_vec_out = 64'b0001111001110101101011101010001011101111100111011001100100101011;
          4:
            level_vec_out = 64'b0001111001110101101011101010001011101111100111011001100100101011;
          5:
            level_vec_out = 64'b1001111001110101101011101010001011101111100111011001100100101011;
          6:
            level_vec_out = 64'b1001111001110101101011101010101011101111100111011001100100101011;
          7:
            level_vec_out = 64'b1001111001110101101111101010101011101111100111011001100100101011;
          8:
            level_vec_out = 64'b1001111001110101101111101010101011101111100111011101100100101011;
          9:
            level_vec_out = 64'b1001111001111101101111101110101011101111100111011101100100101011;
          10:
            level_vec_out = 64'b1011111001111101101111101110101011101111100111011101100100101011;
          11:
            level_vec_out = 64'b1011111001111101101111101110101111101111100111011101100100101011;
          12:
            level_vec_out = 64'b1011111001111101101111101110101111101111100111011101100100101011;
          13:
            level_vec_out = 64'b1011111001111101101111101110101111101111100111011101100101101011;
          14:
            level_vec_out = 64'b1011111011111101101111101111101111101111101111011101100101101011;
          15:
            level_vec_out = 64'b1011111111111101101111101111101111101111101111011111101101101011;
          16:
            level_vec_out = 64'b1011111111111101101111101111101111101111101111111111101101111011;
          17:
            level_vec_out = 64'b1011111111111101101111101111101111101111101111111111101101111011;
          18:
            level_vec_out = 64'b1011111111111111101111101111101111101111101111111111101101111011;
          19:
            level_vec_out = 64'b1011111111111111101111101111111111101111101111111111101101111011;
          20:
            level_vec_out = 64'b1011111111111111101111101111111111101111101111111111101101111011;
          21:
            level_vec_out = 64'b1011111111111111101111101111111111101111101111111111101101111011;
          22:
            level_vec_out = 64'b1011111111111111111111101111111111101111101111111111101101111011;
          23:
            level_vec_out = 64'b1111111111111111111111101111111111101111101111111111101101111011;
          24:
            level_vec_out = 64'b1111111111111111111111101111111111101111101111111111101101111011;
          25:
            level_vec_out = 64'b1111111111111111111111101111111111101111101111111111101101111011;
          26:
            level_vec_out = 64'b1111111111111111111111101111111111101111101111111111101101111011;
          27:
            level_vec_out = 64'b1111111111111111111111101111111111101111111111111111101101111011;
          28:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111101111011;
          29:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111101111011;
          30:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111101111011;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111011;
        endcase
      4:
        case (frame_id)
          0:
            level_vec_out = 64'b1100001000101110111101101011110001000011001001111111011010100000;
          1:
            level_vec_out = 64'b1100001000101110111101101011110001000011001001111111011010100000;
          2:
            level_vec_out = 64'b1100001000101110111111101011110001000011001001111111011010100000;
          3:
            level_vec_out = 64'b1100001000101110111111101011110001000011001001111111011010100000;
          4:
            level_vec_out = 64'b1100001000101110111111101011110011000011001001111111011010100000;
          5:
            level_vec_out = 64'b1100001000101110111111101011110011000011001001111111011010100000;
          6:
            level_vec_out = 64'b1100001000101110111111101011110011000011001001111111011010100000;
          7:
            level_vec_out = 64'b1100001000101110111111101011110011010011001001111111111010100000;
          8:
            level_vec_out = 64'b1100001000101110111111101011110011010011011001111111111010100000;
          9:
            level_vec_out = 64'b1100001000111110111111101011110011010011011001111111111010100000;
          10:
            level_vec_out = 64'b1100001000111110111111101011110011010011011001111111111010100001;
          11:
            level_vec_out = 64'b1100101000111110111111101011110011110011011001111111111010110001;
          12:
            level_vec_out = 64'b1100111000111110111111101011110011111011011001111111111010110001;
          13:
            level_vec_out = 64'b1101111000111110111111101011110011111111011001111111111010110001;
          14:
            level_vec_out = 64'b1101111000111110111111101011110011111111011001111111111010110001;
          15:
            level_vec_out = 64'b1101111001111110111111101011110011111111111001111111111010110001;
          16:
            level_vec_out = 64'b1101111001111110111111101011110011111111111101111111111010110001;
          17:
            level_vec_out = 64'b1101111001111110111111101011110011111111111101111111111010111001;
          18:
            level_vec_out = 64'b1101111011111110111111101011110111111111111101111111111010111001;
          19:
            level_vec_out = 64'b1101111011111110111111101011110111111111111101111111111010111001;
          20:
            level_vec_out = 64'b1101111011111111111111101011111111111111111101111111111010111001;
          21:
            level_vec_out = 64'b1101111011111111111111101011111111111111111101111111111010111001;
          22:
            level_vec_out = 64'b1101111011111111111111101111111111111111111101111111111010111001;
          23:
            level_vec_out = 64'b1101111011111111111111101111111111111111111101111111111010111001;
          24:
            level_vec_out = 64'b1101111011111111111111101111111111111111111101111111111011111001;
          25:
            level_vec_out = 64'b1101111111111111111111101111111111111111111101111111111011111001;
          26:
            level_vec_out = 64'b1101111111111111111111101111111111111111111111111111111111111001;
          27:
            level_vec_out = 64'b1101111111111111111111101111111111111111111111111111111111111011;
          28:
            level_vec_out = 64'b1101111111111111111111111111111111111111111111111111111111111011;
          29:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
          30:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        endcase
      5:
        case (frame_id)
          0:
            level_vec_out = 64'b1001001011101010011001100110101010111010011010100000000011101010;
          1:
            level_vec_out = 64'b1001001011101010011001100110101010111010011010100110000111101010;
          2:
            level_vec_out = 64'b1001001011101010011001100110101010111010011010100110000111101010;
          3:
            level_vec_out = 64'b1001001011101010011001100110101010111010011010101110000111101010;
          4:
            level_vec_out = 64'b1001001011101010011001100110101010111010011010101110000111101110;
          5:
            level_vec_out = 64'b1001001011101010111001100110101010111011011010101110000111101110;
          6:
            level_vec_out = 64'b1001001011111010111001100110101010111011011110101110000111101110;
          7:
            level_vec_out = 64'b1001001011111010111001100110101010111011011110101110000111101110;
          8:
            level_vec_out = 64'b1001001011111010111001100110101010111011011110101110100111101110;
          9:
            level_vec_out = 64'b1001001011111010111001100110101010111011011110101110100111101110;
          10:
            level_vec_out = 64'b1001001011111010111001100110101010111011011110101110100111101110;
          11:
            level_vec_out = 64'b1101001011111010111001100110101010111011011110101110100111101110;
          12:
            level_vec_out = 64'b1101001111111010111001100110101010111011011110101110100111101110;
          13:
            level_vec_out = 64'b1101001111111010111001100111101010111011011110101110100111101110;
          14:
            level_vec_out = 64'b1101001111111010111001100111101010111011011110101110100111101110;
          15:
            level_vec_out = 64'b1101001111111011111001100111101010111011011110101110100111101110;
          16:
            level_vec_out = 64'b1101001111111011111001100111101010111011011110101110100111101110;
          17:
            level_vec_out = 64'b1101001111111011111001100111101010111011011110101110100111101110;
          18:
            level_vec_out = 64'b1101001111111011111001100111101010111011011110101110100111101110;
          19:
            level_vec_out = 64'b1101001111111011111001100111101010111011011110101110100111111110;
          20:
            level_vec_out = 64'b1101001111111111111001100111101010111011011110101110100111111110;
          21:
            level_vec_out = 64'b1101001111111111111001100111101010111011011111101111100111111110;
          22:
            level_vec_out = 64'b1101001111111111111001100111101010111011111111101111100111111110;
          23:
            level_vec_out = 64'b1101001111111111111001111111101010111011111111101111100111111110;
          24:
            level_vec_out = 64'b1101101111111111111001111111101010111111111111101111100111111111;
          25:
            level_vec_out = 64'b1101101111111111111001111111111110111111111111101111100111111111;
          26:
            level_vec_out = 64'b1101101111111111111011111111111110111111111111101111100111111111;
          27:
            level_vec_out = 64'b1101101111111111111111111111111110111111111111101111100111111111;
          28:
            level_vec_out = 64'b1101101111111111111111111111111110111111111111101111100111111111;
          29:
            level_vec_out = 64'b1101101111111111111111111111111110111111111111101111100111111111;
          30:
            level_vec_out = 64'b1111111111111111111111111111111110111111111111111111110111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111110111111111;
        endcase
      6:
        case (frame_id)
          0:
            level_vec_out = 64'b1010010101000011001011100000110101010111011011100110000111010101;
          1:
            level_vec_out = 64'b1010010101000011001011100000110101010111011011100110000111010101;
          2:
            level_vec_out = 64'b1010010101000011001011101000110101010111111011100110000111010101;
          3:
            level_vec_out = 64'b1010010101000011001011101001110101010111111011100110000111010101;
          4:
            level_vec_out = 64'b1010010101000111001011101001111101010111111011100110000111010101;
          5:
            level_vec_out = 64'b1010010101100111001011101001111101010111111011100110001111010101;
          6:
            level_vec_out = 64'b1010010101100111001011101001111101110111111011100110001111010101;
          7:
            level_vec_out = 64'b1010010101100111101011101001111101110111111011100110001111010101;
          8:
            level_vec_out = 64'b1010010101100111101011101101111101110111111011100110011111010101;
          9:
            level_vec_out = 64'b1010010101100111101011101101111101110111111011100110011111010111;
          10:
            level_vec_out = 64'b1010010101100111101011101101111101110111111011100110011111010111;
          11:
            level_vec_out = 64'b1010010111100111101011101101111101110111111011100110011111010111;
          12:
            level_vec_out = 64'b1010010111100111101011101101111101110111111011100110011111010111;
          13:
            level_vec_out = 64'b1010010111100111101011101101111101110111111011100110011111110111;
          14:
            level_vec_out = 64'b1010010111100111101011111101111101110111111011100110011111110111;
          15:
            level_vec_out = 64'b1010010111100111101011111101111101110111111011100110011111110111;
          16:
            level_vec_out = 64'b1010010111100111111011111101111101110111111011100110011111110111;
          17:
            level_vec_out = 64'b1010110111100111111011111101111101110111111011100110011111110111;
          18:
            level_vec_out = 64'b1010110111100111111011111101111101110111111011101110011111110111;
          19:
            level_vec_out = 64'b1010110111100111111011111101111101110111111011101110011111111111;
          20:
            level_vec_out = 64'b1010110111100111111011111101111101110111111111101110011111111111;
          21:
            level_vec_out = 64'b1011110111100111111011111101111101110111111111101110011111111111;
          22:
            level_vec_out = 64'b1011110111100111111011111101111101110111111111111111011111111111;
          23:
            level_vec_out = 64'b1011110111100111111011111101111101111111111111111111111111111111;
          24:
            level_vec_out = 64'b1011111111100111111011111111111101111111111111111111111111111111;
          25:
            level_vec_out = 64'b1011111111100111111011111111111101111111111111111111111111111111;
          26:
            level_vec_out = 64'b1011111111100111111111111111111101111111111111111111111111111111;
          27:
            level_vec_out = 64'b1111111111101111111111111111111101111111111111111111111111111111;
          28:
            level_vec_out = 64'b1111111111101111111111111111111101111111111111111111111111111111;
          29:
            level_vec_out = 64'b1111111111101111111111111111111111111111111111111111111111111111;
          30:
            level_vec_out = 64'b1111111111101111111111111111111111111111111111111111111111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        endcase
      7:
        case (frame_id)
          0:
            level_vec_out = 64'b0101000111001001101111101000000111011010001110100000100001101011;
          1:
            level_vec_out = 64'b0101000111001001101111101000000111011010001110100000100001101011;
          2:
            level_vec_out = 64'b0101000111001001101111101000000111011010001110100000100001101011;
          3:
            level_vec_out = 64'b0101000111001001101111101000100111011011001110100000100001101011;
          4:
            level_vec_out = 64'b0101000111001001101111101100100111011011001110100000100001101011;
          5:
            level_vec_out = 64'b0101000111001001101111101100100111011011001110100010100001101011;
          6:
            level_vec_out = 64'b0101000111011001101111101100100111011011001110100010100001101011;
          7:
            level_vec_out = 64'b0101010111011001101111101100100111011011001110100010100001101111;
          8:
            level_vec_out = 64'b0101010111011001101111101100100111011011001110100010100001101111;
          9:
            level_vec_out = 64'b0101011111011001101111101100100111111011001110100010100001101111;
          10:
            level_vec_out = 64'b0101011111011001111111101100100111111011001111100010100001101111;
          11:
            level_vec_out = 64'b0101011111011001111111101100100111111011001111100010100001101111;
          12:
            level_vec_out = 64'b0101011111011001111111101100100111111011001111100010100001101111;
          13:
            level_vec_out = 64'b0111011111011001111111111100100111111011001111100010100001101111;
          14:
            level_vec_out = 64'b1111011111011001111111111100100111111011001111100010101001101111;
          15:
            level_vec_out = 64'b1111011111011001111111111100100111111011011111100010101001101111;
          16:
            level_vec_out = 64'b1111011111011001111111111101100111111011011111100010101001101111;
          17:
            level_vec_out = 64'b1111011111011101111111111101100111111111011111100010101001101111;
          18:
            level_vec_out = 64'b1111011111011101111111111101100111111111011111100010101001101111;
          19:
            level_vec_out = 64'b1111011111011101111111111101100111111111011111100010101111101111;
          20:
            level_vec_out = 64'b1111011111011101111111111101100111111111011111101111101111101111;
          21:
            level_vec_out = 64'b1111111111011111111111111101100111111111011111101111111111101111;
          22:
            level_vec_out = 64'b1111111111011111111111111111100111111111011111101111111111101111;
          23:
            level_vec_out = 64'b1111111111011111111111111111100111111111011111101111111111101111;
          24:
            level_vec_out = 64'b1111111111011111111111111111100111111111011111101111111111111111;
          25:
            level_vec_out = 64'b1111111111111111111111111111100111111111011111101111111111111111;
          26:
            level_vec_out = 64'b1111111111111111111111111111100111111111011111101111111111111111;
          27:
            level_vec_out = 64'b1111111111111111111111111111100111111111011111101111111111111111;
          28:
            level_vec_out = 64'b1111111111111111111111111111100111111111011111101111111111111111;
          29:
            level_vec_out = 64'b1111111111111111111111111111100111111111011111111111111111111111;
          30:
            level_vec_out = 64'b1111111111111111111111111111110111111111011111111111111111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111110111111111111111111111111111111111;
        endcase
    endcase
  end
endmodule