----
 -- @file level_hvec_gen_hdl.hpp
 -- @brief This script generates HDL code for generating high-dimensional LEVEL vectors.
 -- It is a novel method; for more information, please refer to our paper.
 --
 -- @author Saeid Jamili and Marco Angioli
 -- @note Author names are listed in alphabetical order.
 -- @email <saeid.jamili@uniroma1.it>
 -- @email <marco.angioli@uniroma1.it>
 --
 -- @contributors
 --
 -- @date Created: 24th July 2023
 -- @date Last Updated: 23th August 2023
 --
 -- @version 1.0.0
 --
 -- @institute Sapienza University of Rome
 -- @cite https://doi.org/10.xxxx/yyyyy
 --
 -- @section DEPENDENCIES
 -- - Dependency1: Description or version details.
 -- - Dependency2: Description or version details.
 --
 -- @section LICENSE
 -- This file is part of the Aeneas HyperCompute Platform.
 --
 -- Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 --
 -- @section CHANGELOG
 -- @version 1.0.0-dev - 23th August 2023
 -- - Initial release
 --
 -- @todo
 -- - Complete level vector generator function
 -- - Add training
 --
 -- @see
 -- -
 -- -
 -- -
 --
 --

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity level_vec_gen is
    Port ( level_vec_out : out  STD_LOGIC_VECTOR (63 downto 0);
           frame_index : in  STD_LOGIC_VECTOR (2 downto 0);
           frame_id : in  STD_LOGIC_VECTOR (4 downto 0));
end level_vec_gen;

architecture Behavioral of level_vec_gen is
begin
    process (frame_index, frame_id)
    begin
        -- Update this function to match your requirements
        case frame_index is
            when "000" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0010000110011001001100000000111011001110110010001010010100100010";
                    when "00001" => level_vec_out <= "0010000110011001001100000000111011001110110010001010010100100010";
                    when "00010" => level_vec_out <= "0010000110011001001100010000111011001110110010001010010100100010";
                    when "00011" => level_vec_out <= "0010000110011001001100010000111011001110110010001010010100100010";
                    when "00100" => level_vec_out <= "0010001110011001001100010000111011001110110010001010010100100110";
                    when "00101" => level_vec_out <= "0010001110011001001100010000111011001110110010001011010100100110";
                    when "00110" => level_vec_out <= "1010001110011001001110010000111011001110110010001011010100100110";
                    when "00111" => level_vec_out <= "1010001110011001001110010000111011001110111010001011010100100110";
                    when "01000" => level_vec_out <= "1010001110011001001110010000111011001110111010011011010100100110";
                    when "01001" => level_vec_out <= "1010001110011001011110010000111011001110111010011011010100100110";
                    when "01010" => level_vec_out <= "1010001110011001111111010000111011001110111010011011010100100110";
                    when "01011" => level_vec_out <= "1010001110011001111111010000111011001110111010011011010100100110";
                    when "01100" => level_vec_out <= "1011001110011001111111011000111011001110111010011011010100100110";
                    when "01101" => level_vec_out <= "1011001110011001111111011000111011001110111010011011010100100110";
                    when "01110" => level_vec_out <= "1011001110011001111111011000111011001110111010011011010100100110";
                    when "01111" => level_vec_out <= "1011001110011001111111011000111011001110111010011011010100100110";
                    when "10000" => level_vec_out <= "1011101110011001111111011000111011001110111010011011010100100110";
                    when "10001" => level_vec_out <= "1011101110111001111111011000111011101110111010011011010100100110";
                    when "10010" => level_vec_out <= "1111101110111001111111011000111011101110111010011011010110100110";
                    when "10011" => level_vec_out <= "1111101110111001111111111000111011101110111010011011010110100110";
                    when "10100" => level_vec_out <= "1111111110111001111111111000111011101111111010011011010110100110";
                    when "10101" => level_vec_out <= "1111111111111001111111111000111011111111111010011011010110100111";
                    when "10110" => level_vec_out <= "1111111111111001111111111000111011111111111010011011010110100111";
                    when "10111" => level_vec_out <= "1111111111111001111111111000111011111111111010011011010110101111";
                    when "11000" => level_vec_out <= "1111111111111001111111111010111111111111111010011011010110101111";
                    when "11001" => level_vec_out <= "1111111111111101111111111010111111111111111010011011110110101111";
                    when "11010" => level_vec_out <= "1111111111111101111111111010111111111111111010011011110110101111";
                    when "11011" => level_vec_out <= "1111111111111101111111111010111111111111111111011011110110101111";
                    when "11100" => level_vec_out <= "1111111111111101111111111011111111111111111111011011110110101111";
                    when "11101" => level_vec_out <= "1111111111111101111111111111111111111111111111111011110110101111";
                    when "11110" => level_vec_out <= "1111111111111101111111111111111111111111111111111111110110101111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111110101111";
                when others => null;
                end case;
            when "001" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0111111111110110011111010010111110101111101110010010000110011011";
                    when "00001" => level_vec_out <= "1111111111110110011111010010111110101111101110010010000110011011";
                    when "00010" => level_vec_out <= "1111111111110110111111010010111110101111101110011010100110011011";
                    when "00011" => level_vec_out <= "1111111111110110111111010010111110101111101110011010100110011011";
                    when "00100" => level_vec_out <= "1111111111110110111111010010111110101111101110011010100110011011";
                    when "00101" => level_vec_out <= "1111111111110110111111010010111110101111101110011011100110011111";
                    when "00110" => level_vec_out <= "1111111111110110111111010010111110101111101111011011110110011111";
                    when "00111" => level_vec_out <= "1111111111110110111111010010111110101111101111011011110110011111";
                    when "01000" => level_vec_out <= "1111111111110110111111010010111110101111101111011011110110011111";
                    when "01001" => level_vec_out <= "1111111111110110111111010010111110101111101111011011110110011111";
                    when "01010" => level_vec_out <= "1111111111110110111111010010111110101111101111011011110110011111";
                    when "01011" => level_vec_out <= "1111111111110110111111010010111110101111101111011011110110011111";
                    when "01100" => level_vec_out <= "1111111111110110111111010010111110101111101111011011110110011111";
                    when "01101" => level_vec_out <= "1111111111110110111111010010111110101111101111011011110110011111";
                    when "01110" => level_vec_out <= "1111111111110110111111010010111110101111101111011011111110011111";
                    when "01111" => level_vec_out <= "1111111111110110111111010011111111101111101111011011111110011111";
                    when "10000" => level_vec_out <= "1111111111110110111111010011111111101111101111011011111110011111";
                    when "10001" => level_vec_out <= "1111111111110110111111010011111111111111101111011011111110111111";
                    when "10010" => level_vec_out <= "1111111111110110111111010011111111111111101111011111111110111111";
                    when "10011" => level_vec_out <= "1111111111110110111111110011111111111111101111011111111110111111";
                    when "10100" => level_vec_out <= "1111111111110110111111110011111111111111101111011111111110111111";
                    when "10101" => level_vec_out <= "1111111111110110111111110011111111111111101111011111111110111111";
                    when "10110" => level_vec_out <= "1111111111110110111111110011111111111111101111011111111110111111";
                    when "10111" => level_vec_out <= "1111111111110110111111110011111111111111101111011111111110111111";
                    when "11000" => level_vec_out <= "1111111111110110111111111011111111111111101111011111111110111111";
                    when "11001" => level_vec_out <= "1111111111110111111111111011111111111111101111011111111111111111";
                    when "11010" => level_vec_out <= "1111111111110111111111111011111111111111101111011111111111111111";
                    when "11011" => level_vec_out <= "1111111111110111111111111111111111111111111111011111111111111111";
                    when "11100" => level_vec_out <= "1111111111110111111111111111111111111111111111011111111111111111";
                    when "11101" => level_vec_out <= "1111111111110111111111111111111111111111111111011111111111111111";
                    when "11110" => level_vec_out <= "1111111111110111111111111111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "010" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0011101111100110100010011110100101010101110010100111100001110010";
                    when "00001" => level_vec_out <= "0011101111100110100011011111100111010101110010100111100001110010";
                    when "00010" => level_vec_out <= "0011101111100110100011011111100111010101110010100111100001110010";
                    when "00011" => level_vec_out <= "0011101111101110100011011111100111011101110010100111100001110010";
                    when "00100" => level_vec_out <= "0011101111101110100011011111100111011101110010100111100001110010";
                    when "00101" => level_vec_out <= "0011101111101110100011011111100111011101110010100111100001110010";
                    when "00110" => level_vec_out <= "0011101111101110110011011111100111011101110010100111100001110010";
                    when "00111" => level_vec_out <= "0011101111101110110011011111100111011101110010100111100101110011";
                    when "01000" => level_vec_out <= "0011101111101110110011011111101111011101110010100111110101110011";
                    when "01001" => level_vec_out <= "0011101111101110110011011111101111011101111010100111110101110011";
                    when "01010" => level_vec_out <= "0011101111101110110011111111101111011101111010100111110101110011";
                    when "01011" => level_vec_out <= "0011101111101110110011111111101111011101111011100111110101110011";
                    when "01100" => level_vec_out <= "0011101111101110110011111111111111011101111011100111110101110011";
                    when "01101" => level_vec_out <= "0111101111101110111011111111111111011101111011100111110101110011";
                    when "01110" => level_vec_out <= "0111101111101110111011111111111111011101111011100111110101110011";
                    when "01111" => level_vec_out <= "0111101111101110111011111111111111011101111011100111110101110011";
                    when "10000" => level_vec_out <= "0111101111101111111011111111111111011101111011110111110101110011";
                    when "10001" => level_vec_out <= "0111101111101111111011111111111111011101111011110111110101110011";
                    when "10010" => level_vec_out <= "0111111111101111111011111111111111011101111011110111110101110011";
                    when "10011" => level_vec_out <= "0111111111101111111011111111111111011101111011110111110101110011";
                    when "10100" => level_vec_out <= "0111111111101111111011111111111111011101111011110111110101110011";
                    when "10101" => level_vec_out <= "0111111111101111111011111111111111011101111011110111110101110111";
                    when "10110" => level_vec_out <= "0111111111101111111111111111111111011101111011110111110111110111";
                    when "10111" => level_vec_out <= "1111111111101111111111111111111111011101111111110111110111111111";
                    when "11000" => level_vec_out <= "1111111111101111111111111111111111011101111111110111110111111111";
                    when "11001" => level_vec_out <= "1111111111101111111111111111111111011101111111110111110111111111";
                    when "11010" => level_vec_out <= "1111111111101111111111111111111111011101111111110111110111111111";
                    when "11011" => level_vec_out <= "1111111111101111111111111111111111011101111111110111110111111111";
                    when "11100" => level_vec_out <= "1111111111111111111111111111111111011101111111110111110111111111";
                    when "11101" => level_vec_out <= "1111111111111111111111111111111111011101111111111111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "011" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0001100101101100000010111000011111001000011011110011100100000100";
                    when "00001" => level_vec_out <= "0001100101101100000010111000011111001000011011110011100100000100";
                    when "00010" => level_vec_out <= "0001100101101100000010111000011111001000011011110011100100000100";
                    when "00011" => level_vec_out <= "0001100101101100000010111010011111001000011011110011100100000100";
                    when "00100" => level_vec_out <= "0001100101101100000110111010011111001010011011110011100100000100";
                    when "00101" => level_vec_out <= "0001100101111100000110111010011111101010011011110011100100000100";
                    when "00110" => level_vec_out <= "0001100101111100000110111010011111101010011011110011100100000100";
                    when "00111" => level_vec_out <= "0001100101111110000110111010011111101110111011110011100100000100";
                    when "01000" => level_vec_out <= "0001101101111110000110111010011111111110111011110011100100000100";
                    when "01001" => level_vec_out <= "0011101101111110000110111010011111111110111011110011100100000100";
                    when "01010" => level_vec_out <= "0011101101111110000110111010011111111111111011110011100101000100";
                    when "01011" => level_vec_out <= "0011101101111110000110111010011111111111111011110011100101000100";
                    when "01100" => level_vec_out <= "0011101101111110000110111010011111111111111011110011110101000100";
                    when "01101" => level_vec_out <= "0011101101111110000110111010011111111111111011110011110101000100";
                    when "01110" => level_vec_out <= "0011101101111110000110111110011111111111111011110011110101010100";
                    when "01111" => level_vec_out <= "1011101101111110000110111110111111111111111011110011110101010100";
                    when "10000" => level_vec_out <= "1011101101111110000110111110111111111111111011110011110101010100";
                    when "10001" => level_vec_out <= "1011101101111110000110111110111111111111111011111011110101010101";
                    when "10010" => level_vec_out <= "1011101111111110000110111110111111111111111011111011110101010101";
                    when "10011" => level_vec_out <= "1011101111111110100110111110111111111111111011111111110101010111";
                    when "10100" => level_vec_out <= "1011101111111110100110111110111111111111111011111111111101010111";
                    when "10101" => level_vec_out <= "1011101111111110100110111110111111111111111011111111111101010111";
                    when "10110" => level_vec_out <= "1011101111111110100110111110111111111111111011111111111101010111";
                    when "10111" => level_vec_out <= "1011101111111110101110111110111111111111111011111111111101010111";
                    when "11000" => level_vec_out <= "1011101111111110101110111110111111111111111011111111111101010111";
                    when "11001" => level_vec_out <= "1011101111111110101110111110111111111111111011111111111101010111";
                    when "11010" => level_vec_out <= "1011111111111110101111111110111111111111111011111111111101010111";
                    when "11011" => level_vec_out <= "1011111111111110111111111110111111111111111011111111111101010111";
                    when "11100" => level_vec_out <= "1011111111111110111111111110111111111111111011111111111111010111";
                    when "11101" => level_vec_out <= "1011111111111110111111111110111111111111111011111111111111110111";
                    when "11110" => level_vec_out <= "1011111111111110111111111111111111111111111011111111111111110111";
                    when "11111" => level_vec_out <= "1011111111111110111111111111111111111111111011111111111111111111";
                when others => null;
                end case;
            when "100" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0110010100011010000100010001110011011010101110110011110100001001";
                    when "00001" => level_vec_out <= "0110010100011010000100010001110011011010101110110011110100001001";
                    when "00010" => level_vec_out <= "0110010100011010000100010001110011011010101110110011110100001001";
                    when "00011" => level_vec_out <= "0110010100011010000100010001110011011010101110110011110100001001";
                    when "00100" => level_vec_out <= "0110010110011110000100010001111011011010101110110011110100001001";
                    when "00101" => level_vec_out <= "0110010110011110000100010001111111011010101110110011110100001001";
                    when "00110" => level_vec_out <= "0110010110011110000100010001111111011010101110110011110100001001";
                    when "00111" => level_vec_out <= "0111010110011110000100010001111111011010101110110011110100001001";
                    when "01000" => level_vec_out <= "0111010110011110000100010001111111011110101110110011110100001001";
                    when "01001" => level_vec_out <= "0111010110011110000100010001111111011110111110110011110100001001";
                    when "01010" => level_vec_out <= "0111010110011110000100010001111111011110111110110011110100001001";
                    when "01011" => level_vec_out <= "0111010110011110000100010001111111011110111110110011110100001001";
                    when "01100" => level_vec_out <= "0111010110011110000101010001111111011110111110110011110100001001";
                    when "01101" => level_vec_out <= "0111010110011110000111110001111111011110111110110011110100001001";
                    when "01110" => level_vec_out <= "0111010110011110000111110001111111011110111110110011110110001001";
                    when "01111" => level_vec_out <= "0111010110111110000111110001111111011110111110110011110110001011";
                    when "10000" => level_vec_out <= "0111010110111110010111110011111111011110111111110011110110001011";
                    when "10001" => level_vec_out <= "0111010110111110010111110011111111011110111111110011110110001011";
                    when "10010" => level_vec_out <= "0111010110111110010111110011111111011110111111110011110110001011";
                    when "10011" => level_vec_out <= "0111010110111110010111110011111111011110111111111011110110001011";
                    when "10100" => level_vec_out <= "0111011110111110010111110011111111011110111111111011111110001011";
                    when "10101" => level_vec_out <= "0111111110111110010111110011111111011110111111111011111110001011";
                    when "10110" => level_vec_out <= "0111111111111110110111110111111111011110111111111111111110001111";
                    when "10111" => level_vec_out <= "0111111111111110110111110111111111011110111111111111111110001111";
                    when "11000" => level_vec_out <= "0111111111111110110111110111111111011110111111111111111110001111";
                    when "11001" => level_vec_out <= "0111111111111110111111110111111111011110111111111111111110001111";
                    when "11010" => level_vec_out <= "0111111111111110111111110111111111011110111111111111111110111111";
                    when "11011" => level_vec_out <= "1111111111111110111111110111111111011110111111111111111110111111";
                    when "11100" => level_vec_out <= "1111111111111110111111110111111111011111111111111111111110111111";
                    when "11101" => level_vec_out <= "1111111111111110111111111111111111011111111111111111111110111111";
                    when "11110" => level_vec_out <= "1111111111111110111111111111111111011111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111011111111111111111111111111111";
                when others => null;
                end case;
            when "101" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1101000010011100101101110101110000100010010001101000110011101011";
                    when "00001" => level_vec_out <= "1101000010011100111101110101110000100110010001101000110011101011";
                    when "00010" => level_vec_out <= "1101000011011100111101110101110001110110010001101000110011101011";
                    when "00011" => level_vec_out <= "1101000011011101111101110101110001110110110001101000110011101011";
                    when "00100" => level_vec_out <= "1101000011011101111101110101110001110110110101101000110011101011";
                    when "00101" => level_vec_out <= "1101000011011101111101111101110001110110110101101000110011101011";
                    when "00110" => level_vec_out <= "1101000011011101111101111101110001110110110101101000110011101011";
                    when "00111" => level_vec_out <= "1101000011011101111101111101110001110110110101101000110011101011";
                    when "01000" => level_vec_out <= "1101000011011101111101111101110001110110110101101000110011111011";
                    when "01001" => level_vec_out <= "1101100011011101111101111101110001110110110101101000110011111011";
                    when "01010" => level_vec_out <= "1101100011011101111101111101110001111110110101101000110011111011";
                    when "01011" => level_vec_out <= "1101100011011101111111111101110001111110110101101000110011111011";
                    when "01100" => level_vec_out <= "1101100011011101111111111111110001111110110101101010110011111011";
                    when "01101" => level_vec_out <= "1101100011011101111111111111110001111110110101101010110011111111";
                    when "01110" => level_vec_out <= "1101100011011101111111111111110011111110110101101010110011111111";
                    when "01111" => level_vec_out <= "1101100011011111111111111111110011111110110101101010110011111111";
                    when "10000" => level_vec_out <= "1101100011011111111111111111110011111110110101101010110011111111";
                    when "10001" => level_vec_out <= "1101100011011111111111111111110011111110110101101010110011111111";
                    when "10010" => level_vec_out <= "1101110011011111111111111111110011111110110111101010110011111111";
                    when "10011" => level_vec_out <= "1101110011111111111111111111110011111110110111101010110011111111";
                    when "10100" => level_vec_out <= "1101110011111111111111111111110011111110110111101010110011111111";
                    when "10101" => level_vec_out <= "1101110011111111111111111111110011111110110111101110110011111111";
                    when "10110" => level_vec_out <= "1101110011111111111111111111110011111110110111101110110011111111";
                    when "10111" => level_vec_out <= "1101110011111111111111111111110011111110111111101110110011111111";
                    when "11000" => level_vec_out <= "1101110011111111111111111111110111111111111111101111110011111111";
                    when "11001" => level_vec_out <= "1101110011111111111111111111110111111111111111101111110111111111";
                    when "11010" => level_vec_out <= "1101110011111111111111111111111111111111111111101111110111111111";
                    when "11011" => level_vec_out <= "1101110011111111111111111111111111111111111111101111110111111111";
                    when "11100" => level_vec_out <= "1111110011111111111111111111111111111111111111101111110111111111";
                    when "11101" => level_vec_out <= "1111110011111111111111111111111111111111111111111111110111111111";
                    when "11110" => level_vec_out <= "1111111011111111111111111111111111111111111111111111110111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111110111111111";
                when others => null;
                end case;
            when "110" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0110101001111100110011101011100111001010011001011100001001010000";
                    when "00001" => level_vec_out <= "0110101001111100110011101011100111011010011001011100001001010000";
                    when "00010" => level_vec_out <= "0110101011111100110011101011100111011010011001011100001001010000";
                    when "00011" => level_vec_out <= "0110101011111110110011101011100111011010011001011100001001010000";
                    when "00100" => level_vec_out <= "0110101011111110110011101011100111011010011001011100001001010000";
                    when "00101" => level_vec_out <= "0110101011111110110011101011100111011010011001011100001001010000";
                    when "00110" => level_vec_out <= "0110101011111110110011101011100111011010011001111100001001010100";
                    when "00111" => level_vec_out <= "0110101011111110110011101011100111011010011001111100001001010100";
                    when "01000" => level_vec_out <= "0110101011111110110011101011100111011010011001111100001001010100";
                    when "01001" => level_vec_out <= "0110101011111110110011101011101111011110011001111100001001010100";
                    when "01010" => level_vec_out <= "0110101011111110110011101011101111011110011001111100001001010100";
                    when "01011" => level_vec_out <= "0110111011111110110011101011101111011110011001111100101011010100";
                    when "01100" => level_vec_out <= "0110111011111110110011101011101111011110011001111100101011010100";
                    when "01101" => level_vec_out <= "0110111011111110110011111011101111111110011001111100101011010100";
                    when "01110" => level_vec_out <= "0110111011111110110011111011101111111110011001111100101111010100";
                    when "01111" => level_vec_out <= "0110111011111110110011111011101111111110011001111100101111010101";
                    when "10000" => level_vec_out <= "0110111011111110111011111011101111111110011001111100101111010101";
                    when "10001" => level_vec_out <= "0110111011111110111011111011101111111110111001111101101111010101";
                    when "10010" => level_vec_out <= "0110111011111110111011111011101111111110111001111101101111010101";
                    when "10011" => level_vec_out <= "0110111011111110111011111011101111111110111001111101101111010101";
                    when "10100" => level_vec_out <= "0110111011111110111011111011101111111110111001111101101111010101";
                    when "10101" => level_vec_out <= "0110111011111110111111111011101111111110111001111101101111010101";
                    when "10110" => level_vec_out <= "0110111011111110111111111011111111111110111001111101101111010101";
                    when "10111" => level_vec_out <= "0110111011111110111111111011111111111110111001111101101111010111";
                    when "11000" => level_vec_out <= "0110111011111110111111111011111111111110111101111101101111010111";
                    when "11001" => level_vec_out <= "0110111011111110111111111011111111111110111101111111101111010111";
                    when "11010" => level_vec_out <= "0110111111111110111111111011111111111110111111111111101111010111";
                    when "11011" => level_vec_out <= "0110111111111110111111111011111111111110111111111111101111110111";
                    when "11100" => level_vec_out <= "1110111111111110111111111111111111111110111111111111111111110111";
                    when "11101" => level_vec_out <= "1110111111111110111111111111111111111110111111111111111111111111";
                    when "11110" => level_vec_out <= "1110111111111111111111111111111111111110111111111111111111111111";
                    when "11111" => level_vec_out <= "1110111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "111" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0011100110010111000111100100010100011101010100111001011110110101";
                    when "00001" => level_vec_out <= "0011100110010111000111100100010100011101010100111001011110111101";
                    when "00010" => level_vec_out <= "0011100110010111000111100100010100011101010100111001011110111101";
                    when "00011" => level_vec_out <= "0011100110010111000111100100010100011101010100111011011111111101";
                    when "00100" => level_vec_out <= "0011100110010111000111100100010100011101010100111011011111111101";
                    when "00101" => level_vec_out <= "1011100110010111000111100100010100011101010100111011011111111101";
                    when "00110" => level_vec_out <= "1011100110010111000111100100010110011101010100111011011111111101";
                    when "00111" => level_vec_out <= "1011100110010111000111100100010110011101010110111011011111111101";
                    when "01000" => level_vec_out <= "1011100110010111000111100100010110011101010110111111011111111101";
                    when "01001" => level_vec_out <= "1011100110010111000111100100010110011101010111111111011111111101";
                    when "01010" => level_vec_out <= "1011100110010111100111100100010110011101010111111111011111111111";
                    when "01011" => level_vec_out <= "1011111110010111100111101100010110011101010111111111011111111111";
                    when "01100" => level_vec_out <= "1011111110010111100111101100110110011101010111111111011111111111";
                    when "01101" => level_vec_out <= "1011111110010111100111101101110110011101010111111111011111111111";
                    when "01110" => level_vec_out <= "1011111110010111100111101101111110011101011111111111011111111111";
                    when "01111" => level_vec_out <= "1011111110010111100111101101111110011101011111111111011111111111";
                    when "10000" => level_vec_out <= "1011111110011111100111101101111110011101011111111111011111111111";
                    when "10001" => level_vec_out <= "1011111110011111100111101101111110011101011111111111011111111111";
                    when "10010" => level_vec_out <= "1011111111011111100111101101111110011101011111111111011111111111";
                    when "10011" => level_vec_out <= "1011111111011111101111101101111110011101011111111111011111111111";
                    when "10100" => level_vec_out <= "1011111111011111111111101111111110011111011111111111011111111111";
                    when "10101" => level_vec_out <= "1011111111011111111111101111111110011111011111111111111111111111";
                    when "10110" => level_vec_out <= "1011111111011111111111101111111110011111011111111111111111111111";
                    when "10111" => level_vec_out <= "1011111111011111111111101111111110111111011111111111111111111111";
                    when "11000" => level_vec_out <= "1111111111011111111111101111111110111111011111111111111111111111";
                    when "11001" => level_vec_out <= "1111111111011111111111101111111111111111011111111111111111111111";
                    when "11010" => level_vec_out <= "1111111111011111111111101111111111111111111111111111111111111111";
                    when "11011" => level_vec_out <= "1111111111111111111111101111111111111111111111111111111111111111";
                    when "11100" => level_vec_out <= "1111111111111111111111101111111111111111111111111111111111111111";
                    when "11101" => level_vec_out <= "1111111111111111111111101111111111111111111111111111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111101111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when others => null;
        end case;
    end process;
end Behavioral;