
/**
 * @file class_hvec_gen_hdl.hpp
 * @brief This script generates HDL code for generating high-dimensional class vectors.
 * It is a novel method; for more information, please refer to our paper.
 *
 * @author Saeid Jamili and Marco Angioli
 * @note Author names are listed in alphabetical order.
 * @email <saeid.jamili@uniroma1.it>
 * @email <marco.angioli@uniroma1.it>
 *
 * @contributors
 *
 * @date Created: 24th July 2023
 * @date Last Updated: 23th August 2023
 *
 * @version 1.0.0
 *
 * @institute Sapienza University of Rome
 * @cite https://doi.org/10.xxxx/yyyyy
 *
 * @section DEPENDENCIES
 * - Dependency1: Description or version details.
 * - Dependency2: Description or version details.
 *
 * @section LICENSE
 * This file is part of the Aeneas HyperCompute Platform.
 *
 * Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 *
 * @section CHANGELOG
 * @version 1.0.0-dev - 23th August 2023
 * - Initial release
 *
 * @todo
 * - Complete level vector generator function
 * - Add training
 *
 * @see
 * -
 * -
 * -
 *
 */

module class_hvec_gen #(parameter int DI_PARALLEL_W_BITS = 64) (
  input logic [2:0] frame_id,
  input logic [1:0] frame_index,
  output logic [DI_PARALLEL_W_BITS-1:0] class_vec_out
);
  always_comb begin
    case (frame_id)
      0:
        case (frame_index)
          0:
            class_vec_out = 64'b371245124521812451224124501094124512452580124501243101601194264012454411228012450124511600115889811381073727612450124570998767124512452312451312451245124571827147181245124510912450001245;
          1:
            class_vec_out = 64'b332232231362232102230167223223300223022120901731102235122102230223199015616614710117342230223211983322322317223402232232231723451082232237223000223;
          2:
            class_vec_out = 64'b91261264112612312609412612680126012399010124012697121012601268801041091050082271260126593810141261262512628126126126733739212612635126000126;
        endcase
      1:
        case (frame_index)
          0:
            class_vec_out = 64'b06600124501245213124514812451245124554701830124512261245538124401541245124512453800124512182941245122624712391245504124512452061348841245177141245015501531094123401041245124500651124572560796;
          1:
            class_vec_out = 64'b018802230223922392232232231840502232142231472230472232232239602232176822322030222223107223223637157223943223095030207222052232230017922310000107;
          2:
            class_vec_out = 64'b168012601266312616126126126570140126124126991160511261261267501261233112612322124126451231261252651267519126082042841260361261260063126810020;
        endcase
      2:
        case (frame_index)
          0:
            class_vec_out = 64'b15268201245700074621245716124590310001044123801222010571245008130500124511561245678618123505280012381245103931236124518300411245698585000123911385381245124501078001245;
          1:
            class_vec_out = 64'b14110602230000770223101223205202158219020801822230019308222312522319363222013100213223001902152233300722316117200021221073223223021400223;
          2:
            class_vec_out = 64'b34710126200051012687126958954123011208612600670261267912668421260480012112600521251264500412695950001208482126126010900126;
        endcase
      3:
        case (frame_index)
          0:
            class_vec_out = 64'b1196066124512201245112212458860002001245751196159103220819280009550001141245012451245169012451245012450119012451223123912456811245124501243495001245016701245124502151074;
          1:
            class_vec_out = 64'b17502223196223101223188000138223822160215101021000097000622302232239502232230223031223220221223197223223022388002230660223223071142;
          2:
            class_vec_out = 64'b1140181261181264412636000531261510578160188800081000311260126126410126126012604441261221261269112612601212300126025012612607071;
        endcase
      4:
        case (frame_index)
          0:
            class_vec_out = 64'b94124512451245108912436941206124510124585012451771245173812451245001245124512459963601245120601364052400058412451019239124501998061166670124550678712451245012451239124557401245019655401245515;
          1:
            class_vec_out = 64'b12232232232072221301902234922314722320223171022322300223223223216902232180338128000105223826223031831782112231021732232230223216223910223018614022377;
          2:
            class_vec_out = 64'b51261261269912697104126291268912649126500126126001261261264816012610104523610008712674221260106270981263371126126012612012647012606795612621;
        endcase
      5:
        case (frame_index)
          0:
            class_vec_out = 64'b903803120473124500641825624012451245012451439901245310008880103012530212451204440612453201245124212451218001200114512450124592504029315400406214012451245625001245280;
          1:
            class_vec_out = 64'b119301640862230029994912223223022315002233200870212173522322339162231922322322321600220219223022369903421001033462232231130022340;
          2:
            class_vec_out = 64'b2413034043126003327715126126012604601260007301094134126125641512637126110126960012464126012625370734100250411261267200126130;
        endcase
      6:
        case (frame_index)
          0:
            class_vec_out = 64'b0105410011245987540114512451245070578663947508052212451245124512451243005777400144124501245321245014307363686110001131232350543029290006880834108802959410121401231;
          1:
            class_vec_out = 64'b0771872231335022122322300014581139124014222322322322322200201166013223022328223091020451650005122325400441700460203214011020501960222;
          2:
            class_vec_out = 64'b095102126752011012612601204378459908112612612612610900564607512601261912603807944310007116456026800073011410706010001230126;
        endcase
      7:
        case (frame_index)
          0:
            class_vec_out = 64'b12450124512450663831245124560912450122600053201245124512451216979312451098010970123612451245012141245124501245124212451245131245246124508671245124568201119124504461245012311374900124501245;
          1:
            class_vec_out = 64'b22302232230420522322377223021300055022322322319721812231580219022122322302132232230223223223223322359223021322322317607222301582230213764502230223;
          2:
            class_vec_out = 64'b12601261260266212612683126012100034012612612610462412611309701261261260122126126012612212612614126601260104126126960451260551260121553201260126;
        endcase
    endcase
  end
endmodule