/**
 * @file level_hvec_gen_hdl.hpp
 * @brief This script generates HDL code for generating high-dimensional LEVEL vectors.
 * It is a novel method; for more information, please refer to our paper.
 *
 * @author Saeid Jamili and Marco Angioli
 * @note Author names are listed in alphabetical order.
 * @email <saeid.jamili@uniroma1.it>
 * @email <marco.angioli@uniroma1.it>
 *
 * @contributors
 *
 * @date Created: 24th July 2023
 * @date Last Updated: 23th August 2023
 *
 * @version 1.0.0
 *
 * @institute Sapienza University of Rome
 * @cite https://doi.org/10.xxxx/yyyyy
 *
 * @section DEPENDENCIES
 * - Dependency1: Description or version details.
 * - Dependency2: Description or version details.
 *
 * @section LICENSE
 * This file is part of the Aeneas HyperCompute Platform.
 *
 * Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 *
 * @section CHANGELOG
 * @version 1.0.0-dev - 23th August 2023
 * - Initial release
 *
 * @todo
 * - Complete level vector generator function
 * - Add training
 *
 * @see
 * -
 * -
 * -
 *
 */

module level_hvec_gen #(parameter int DI_PARALLEL_W_BITS = 64) (
  input logic [2:0] frame_index,
  input logic [4:0] frame_id,
  output logic [DI_PARALLEL_W_BITS-1:0] level_vec_out
);
  always_comb begin
    case (frame_index)
      0:
        case (frame_id)
          0:
            level_vec_out = 64'b1000110001000110010100111010011110011001100111101100001011111001;
          1:
            level_vec_out = 64'b1000110001000110010100111010011110011001100111101100001011111001;
          2:
            level_vec_out = 64'b1000110001000110010100111010011110011001100111101100001011111001;
          3:
            level_vec_out = 64'b1000110001000110010100111010011110011001100111101100001011111001;
          4:
            level_vec_out = 64'b1000110001000110010100111011011110011001100111101100001011111001;
          5:
            level_vec_out = 64'b1000110001010110010100111011011110011101100111101100001011111001;
          6:
            level_vec_out = 64'b1000110001010110010100111011011110011101100111101100011011111001;
          7:
            level_vec_out = 64'b1000110001010110010100111011011110111101100111101100011011111011;
          8:
            level_vec_out = 64'b1000110101010110010100111011011110111101100111101100011011111011;
          9:
            level_vec_out = 64'b1000110101010110010100111011011110111101100111101100011011111011;
          10:
            level_vec_out = 64'b1000110101010110010100111011011110111101100111101100011011111011;
          11:
            level_vec_out = 64'b1000110101010110010100111011011110111101100111101100011011111011;
          12:
            level_vec_out = 64'b1000110101010110011100111011011110111101110111101110011011111111;
          13:
            level_vec_out = 64'b1000110101011110011100111011011110111101110111101110011011111111;
          14:
            level_vec_out = 64'b1000110101011110011100111011011110111101110111101110011011111111;
          15:
            level_vec_out = 64'b1000110101011110011100111011011110111101110111101110011011111111;
          16:
            level_vec_out = 64'b1100110101011110011100111011011110111101110111111110011011111111;
          17:
            level_vec_out = 64'b1100110101011110011100111011011111111101110111111110011011111111;
          18:
            level_vec_out = 64'b1100110101011111011100111011011111111111110111111110011011111111;
          19:
            level_vec_out = 64'b1100110101011111011100111011011111111111110111111111011011111111;
          20:
            level_vec_out = 64'b1100110101111111011100111011011111111111110111111111011011111111;
          21:
            level_vec_out = 64'b1100110101111111011100111011011111111111110111111111011011111111;
          22:
            level_vec_out = 64'b1100110101111111011101111111011111111111110111111111111011111111;
          23:
            level_vec_out = 64'b1100110101111111011101111111011111111111111111111111111011111111;
          24:
            level_vec_out = 64'b1100110101111111011101111111011111111111111111111111111011111111;
          25:
            level_vec_out = 64'b1100110101111111111101111111011111111111111111111111111111111111;
          26:
            level_vec_out = 64'b1100111101111111111101111111011111111111111111111111111111111111;
          27:
            level_vec_out = 64'b1100111101111111111101111111111111111111111111111111111111111111;
          28:
            level_vec_out = 64'b1100111111111111111101111111111111111111111111111111111111111111;
          29:
            level_vec_out = 64'b1100111111111111111101111111111111111111111111111111111111111111;
          30:
            level_vec_out = 64'b1101111111111111111111111111111111111111111111111111111111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        endcase
      1:
        case (frame_id)
          0:
            level_vec_out = 64'b1010001010001000110101011111110010110010101001111010110111010101;
          1:
            level_vec_out = 64'b1010001010001001110101011111111010110010101001111010110111010101;
          2:
            level_vec_out = 64'b1010001010001001110101011111111010110010101001111010111111010101;
          3:
            level_vec_out = 64'b1010001010001001110101011111111010110010101001111010111111010101;
          4:
            level_vec_out = 64'b1010001010001001110101011111111010110010111001111010111111010111;
          5:
            level_vec_out = 64'b1010001010001001110101011111111010110010111001111010111111010111;
          6:
            level_vec_out = 64'b1010001010001001110101011111111010110010111001111010111111010111;
          7:
            level_vec_out = 64'b1010001010011001110101011111111010110010111001111010111111010111;
          8:
            level_vec_out = 64'b1010001010011001110101011111111010110010111001111010111111010111;
          9:
            level_vec_out = 64'b1010011010011001110101011111111010110010111001111010111111010111;
          10:
            level_vec_out = 64'b1010011010011001110101011111111010110010111001111010111111110111;
          11:
            level_vec_out = 64'b1010011010011001110101011111111010110010111001111010111111110111;
          12:
            level_vec_out = 64'b1010011011011001110101011111111010110010111001111010111111110111;
          13:
            level_vec_out = 64'b1110011011011001110101011111111010110010111001111011111111110111;
          14:
            level_vec_out = 64'b1110011011011001110101011111111010110010111001111011111111110111;
          15:
            level_vec_out = 64'b1110111011011001111101011111111010110010111001111011111111111111;
          16:
            level_vec_out = 64'b1110111111011001111101011111111010110110111001111011111111111111;
          17:
            level_vec_out = 64'b1110111111011001111101011111111010110110111001111011111111111111;
          18:
            level_vec_out = 64'b1110111111011001111101011111111010110110111001111011111111111111;
          19:
            level_vec_out = 64'b1110111111011001111101011111111010110110111001111011111111111111;
          20:
            level_vec_out = 64'b1111111111011001111101011111111010110110111001111011111111111111;
          21:
            level_vec_out = 64'b1111111111111001111101011111111110110110111001111011111111111111;
          22:
            level_vec_out = 64'b1111111111111001111101011111111111110110111101111011111111111111;
          23:
            level_vec_out = 64'b1111111111111001111101011111111111110110111101111011111111111111;
          24:
            level_vec_out = 64'b1111111111111001111101111111111111110110111111111011111111111111;
          25:
            level_vec_out = 64'b1111111111111001111101111111111111111110111111111011111111111111;
          26:
            level_vec_out = 64'b1111111111111001111101111111111111111110111111111011111111111111;
          27:
            level_vec_out = 64'b1111111111111001111101111111111111111110111111111011111111111111;
          28:
            level_vec_out = 64'b1111111111111001111111111111111111111111111111111011111111111111;
          29:
            level_vec_out = 64'b1111111111111001111111111111111111111111111111111111111111111111;
          30:
            level_vec_out = 64'b1111111111111001111111111111111111111111111111111111111111111111;
          31:
            level_vec_out = 64'b1111111111111011111111111111111111111111111111111111111111111111;
        endcase
      2:
        case (frame_id)
          0:
            level_vec_out = 64'b0111001110010010101110110001111011011101111011011111100001111011;
          1:
            level_vec_out = 64'b1111001110010010101110110001111011011101111011011111100001111011;
          2:
            level_vec_out = 64'b1111001110010010101110110001111011011101111011011111100101111011;
          3:
            level_vec_out = 64'b1111001110010010101110110001111011011101111111011111100101111011;
          4:
            level_vec_out = 64'b1111001110010010101110110001111011011101111111011111100101111011;
          5:
            level_vec_out = 64'b1111001110010010101110110001111011011111111111011111100101111011;
          6:
            level_vec_out = 64'b1111001110010010101110110001111011011111111111011111100101111011;
          7:
            level_vec_out = 64'b1111001110010010101110110001111011011111111111011111100101111011;
          8:
            level_vec_out = 64'b1111001110110010101110110011111011011111111111011111100101111011;
          9:
            level_vec_out = 64'b1111001110110010101110110011111011011111111111011111110101111011;
          10:
            level_vec_out = 64'b1111001110110010111110111011111011011111111111011111111101111011;
          11:
            level_vec_out = 64'b1111001110110010111110111011111011111111111111011111111101111011;
          12:
            level_vec_out = 64'b1111001110110010111110111011111011111111111111011111111101111011;
          13:
            level_vec_out = 64'b1111001110110010111110111011111011111111111111011111111101111011;
          14:
            level_vec_out = 64'b1111001110110010111110111011111011111111111111011111111101111011;
          15:
            level_vec_out = 64'b1111001110110010111110111011111011111111111111011111111101111011;
          16:
            level_vec_out = 64'b1111001110110010111110111011111011111111111111011111111101111011;
          17:
            level_vec_out = 64'b1111001110110010111111111011111011111111111111011111111101111011;
          18:
            level_vec_out = 64'b1111001110110010111111111011111011111111111111011111111101111011;
          19:
            level_vec_out = 64'b1111001110110010111111111011111011111111111111011111111101111011;
          20:
            level_vec_out = 64'b1111001110110010111111111011111011111111111111011111111101111111;
          21:
            level_vec_out = 64'b1111001110110011111111111011111011111111111111111111111101111111;
          22:
            level_vec_out = 64'b1111001110110011111111111011111011111111111111111111111101111111;
          23:
            level_vec_out = 64'b1111001110110011111111111011111111111111111111111111111101111111;
          24:
            level_vec_out = 64'b1111001111110111111111111011111111111111111111111111111101111111;
          25:
            level_vec_out = 64'b1111101111111111111111111011111111111111111111111111111101111111;
          26:
            level_vec_out = 64'b1111101111111111111111111011111111111111111111111111111101111111;
          27:
            level_vec_out = 64'b1111101111111111111111111011111111111111111111111111111101111111;
          28:
            level_vec_out = 64'b1111101111111111111111111111111111111111111111111111111101111111;
          29:
            level_vec_out = 64'b1111101111111111111111111111111111111111111111111111111101111111;
          30:
            level_vec_out = 64'b1111101111111111111111111111111111111111111111111111111111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        endcase
      3:
        case (frame_id)
          0:
            level_vec_out = 64'b0111111001001100111101100100000010111010000100011001011100011001;
          1:
            level_vec_out = 64'b0111111001001100111101100100000010111010000100011001011100011001;
          2:
            level_vec_out = 64'b0111111001001100111101100100000010111010010100011001011100011001;
          3:
            level_vec_out = 64'b0111111001101100111101100100000010111010111100011001011100011101;
          4:
            level_vec_out = 64'b0111111001101100111101100100000010111010111100011001011110011101;
          5:
            level_vec_out = 64'b0111111001101100111101100100000010111010111100011001111110011101;
          6:
            level_vec_out = 64'b0111111011101100111101101100000010111010111100011001111111011101;
          7:
            level_vec_out = 64'b0111111011101100111101101100000010111010111100011001111111111101;
          8:
            level_vec_out = 64'b0111111011101100111101101100000010111010111110111001111111111101;
          9:
            level_vec_out = 64'b0111111011101100111101101110000010111010111110111001111111111101;
          10:
            level_vec_out = 64'b0111111011101100111101101110000010111010111110111001111111111101;
          11:
            level_vec_out = 64'b0111111011101100111101101110000010111010111110111001111111111101;
          12:
            level_vec_out = 64'b0111111011101100111101101110000010111010111110111011111111111101;
          13:
            level_vec_out = 64'b0111111011101100111101101110000010111010111110111011111111111101;
          14:
            level_vec_out = 64'b0111111011101100111101101110100010111010111110111011111111111101;
          15:
            level_vec_out = 64'b0111111011101100111101101110100010111010111110111011111111111101;
          16:
            level_vec_out = 64'b0111111011101100111101101110100010111010111110111011111111111101;
          17:
            level_vec_out = 64'b0111111111101100111111101110100010111010111110111011111111111101;
          18:
            level_vec_out = 64'b0111111111111100111111101110100110111010111111111011111111111101;
          19:
            level_vec_out = 64'b0111111111111110111111101110100110111010111111111011111111111101;
          20:
            level_vec_out = 64'b0111111111111110111111101110100110111010111111111011111111111101;
          21:
            level_vec_out = 64'b0111111111111110111111101110100110111110111111111011111111111101;
          22:
            level_vec_out = 64'b0111111111111110111111101110100110111110111111111011111111111111;
          23:
            level_vec_out = 64'b1111111111111110111111101110100110111110111111111011111111111111;
          24:
            level_vec_out = 64'b1111111111111110111111101110101110111110111111111011111111111111;
          25:
            level_vec_out = 64'b1111111111111110111111101110101110111110111111111011111111111111;
          26:
            level_vec_out = 64'b1111111111111110111111101110101110111110111111111111111111111111;
          27:
            level_vec_out = 64'b1111111111111110111111101110101110111110111111111111111111111111;
          28:
            level_vec_out = 64'b1111111111111111111111111110101110111110111111111111111111111111;
          29:
            level_vec_out = 64'b1111111111111111111111111110101111111110111111111111111111111111;
          30:
            level_vec_out = 64'b1111111111111111111111111110101111111110111111111111111111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111110101111111111111111111111111111111111;
        endcase
      4:
        case (frame_id)
          0:
            level_vec_out = 64'b0101000001111110110001011000111001010111110010010001100100101000;
          1:
            level_vec_out = 64'b0101000001111110110101011010111001010111110010011001100100101000;
          2:
            level_vec_out = 64'b0101000001111110110101011010111001010111110010011001100100101001;
          3:
            level_vec_out = 64'b0101000001111110110101011010111001010111111010011001100100101001;
          4:
            level_vec_out = 64'b0101000001111110110101011010111001010111111111011001100100101001;
          5:
            level_vec_out = 64'b0101000001111110110101011011111011010111111111011001100100101001;
          6:
            level_vec_out = 64'b0101000001111110110101011011111011010111111111011001100100101001;
          7:
            level_vec_out = 64'b0101000001111110110101011011111011010111111111111001100100101001;
          8:
            level_vec_out = 64'b0101000001111110110101011011111011010111111111111001100100101001;
          9:
            level_vec_out = 64'b0101000001111110110101011011111011010111111111111001110100101001;
          10:
            level_vec_out = 64'b0101000001111110110101011011111111010111111111111001110100101011;
          11:
            level_vec_out = 64'b0101000001111110110101011011111111010111111111111011110100101011;
          12:
            level_vec_out = 64'b0101000001111110110101011011111111010111111111111011110100101011;
          13:
            level_vec_out = 64'b0101000001111110110101011011111111010111111111111011110110101011;
          14:
            level_vec_out = 64'b0101010001111110110111011011111111011111111111111011110110101011;
          15:
            level_vec_out = 64'b0101010001111110110111011111111111011111111111111011110110101011;
          16:
            level_vec_out = 64'b0101010101111110110111011111111111011111111111111011110110101011;
          17:
            level_vec_out = 64'b0101010101111110110111011111111111111111111111111011110110111011;
          18:
            level_vec_out = 64'b0101010101111110110111011111111111111111111111111011110110111011;
          19:
            level_vec_out = 64'b0101010101111110110111011111111111111111111111111011111110111011;
          20:
            level_vec_out = 64'b0101010101111110110111011111111111111111111111111011111110111011;
          21:
            level_vec_out = 64'b0101010101111110110111011111111111111111111111111011111110111011;
          22:
            level_vec_out = 64'b0101010101111110110111011111111111111111111111111011111110111111;
          23:
            level_vec_out = 64'b0101011101111110110111011111111111111111111111111011111110111111;
          24:
            level_vec_out = 64'b0101011101111110110111011111111111111111111111111011111110111111;
          25:
            level_vec_out = 64'b0101011101111110110111011111111111111111111111111011111110111111;
          26:
            level_vec_out = 64'b0101011101111111110111011111111111111111111111111011111110111111;
          27:
            level_vec_out = 64'b1111011101111111111111111111111111111111111111111011111110111111;
          28:
            level_vec_out = 64'b1111111101111111111111111111111111111111111111111011111110111111;
          29:
            level_vec_out = 64'b1111111101111111111111111111111111111111111111111011111110111111;
          30:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111110111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111110111111;
        endcase
      5:
        case (frame_id)
          0:
            level_vec_out = 64'b1101100000010001101011001001110101000111010001100110101110010010;
          1:
            level_vec_out = 64'b1101100000010001101011001001110101000111010001100110101110010010;
          2:
            level_vec_out = 64'b1101100000010011101011101001111101000111010001100110101110010010;
          3:
            level_vec_out = 64'b1101100000010011101011101001111101000111010001110110101110010010;
          4:
            level_vec_out = 64'b1101100000010011101011101001111101000111010001110110101110010010;
          5:
            level_vec_out = 64'b1101100000010011101011101001111101000111010001110110101110010010;
          6:
            level_vec_out = 64'b1101100000010011101011101001111101000111010001110111101110010010;
          7:
            level_vec_out = 64'b1101100000010111101011101001111101000111010001110111101110010010;
          8:
            level_vec_out = 64'b1101100000010111101011101001111101000111010001110111111110010010;
          9:
            level_vec_out = 64'b1101100000010111101011101001111101000111010001110111111110010011;
          10:
            level_vec_out = 64'b1101100000010111101011101001111101000111010001110111111110010011;
          11:
            level_vec_out = 64'b1101100000010111101011101001111101000111110001111111111110010011;
          12:
            level_vec_out = 64'b1101100000010111101011101001111101000111110001111111111110010111;
          13:
            level_vec_out = 64'b1101100000011111101011101001111101000111111001111111111110010111;
          14:
            level_vec_out = 64'b1101110000011111101111101001111101010111111001111111111110010111;
          15:
            level_vec_out = 64'b1101110100011111101111101001111101011111111001111111111110010111;
          16:
            level_vec_out = 64'b1101110100011111101111101001111101011111111001111111111110110111;
          17:
            level_vec_out = 64'b1101110100011111101111101001111101011111111001111111111110110111;
          18:
            level_vec_out = 64'b1101110100011111101111101001111101011111111001111111111110110111;
          19:
            level_vec_out = 64'b1101110100011111101111101001111101111111111001111111111111110111;
          20:
            level_vec_out = 64'b1101110100011111101111101001111101111111111001111111111111110111;
          21:
            level_vec_out = 64'b1101110100011111101111101001111101111111111001111111111111110111;
          22:
            level_vec_out = 64'b1101110100011111101111101001111101111111111001111111111111110111;
          23:
            level_vec_out = 64'b1101110110011111101111101001111101111111111001111111111111110111;
          24:
            level_vec_out = 64'b1101110110011111101111101101111111111111111011111111111111110111;
          25:
            level_vec_out = 64'b1101110110111111111111101101111111111111111011111111111111110111;
          26:
            level_vec_out = 64'b1101110111111111111111101101111111111111111011111111111111110111;
          27:
            level_vec_out = 64'b1111110111111111111111101101111111111111111011111111111111110111;
          28:
            level_vec_out = 64'b1111110111111111111111111101111111111111111011111111111111110111;
          29:
            level_vec_out = 64'b1111111111111111111111111101111111111111111011111111111111111111;
          30:
            level_vec_out = 64'b1111111111111111111111111111111111111111111011111111111111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111011111111111111111111;
        endcase
      6:
        case (frame_id)
          0:
            level_vec_out = 64'b0100010101100101110000010010011010011000100100111110101100001111;
          1:
            level_vec_out = 64'b0100010101100101110000010010011010011000101100111110101100001111;
          2:
            level_vec_out = 64'b0100010101100101110000010010011010011000101101111110101100001111;
          3:
            level_vec_out = 64'b0100010101110101110000010010011010011000101101111110101100001111;
          4:
            level_vec_out = 64'b0100011101110101110000110010011010011000101101111110101100001111;
          5:
            level_vec_out = 64'b0100011101110101110000110010011010011000101101111110101100001111;
          6:
            level_vec_out = 64'b0100011101110101110000110010011010011000101101111110101100001111;
          7:
            level_vec_out = 64'b0100011101110101110010110010011010011000101101111110101100101111;
          8:
            level_vec_out = 64'b0100011101110101110010110010011011011000101101111110101100101111;
          9:
            level_vec_out = 64'b0100011101110101110010110110011011011000101101111110101100101111;
          10:
            level_vec_out = 64'b0100011101110101110010110111011011011000101101111110101110101111;
          11:
            level_vec_out = 64'b0100011111110101110011110111011011011000101101111110101110101111;
          12:
            level_vec_out = 64'b0100011111110101110011110111011011011000101101111110101110101111;
          13:
            level_vec_out = 64'b0100011111110101110011110111011011011000101101111110101110101111;
          14:
            level_vec_out = 64'b0100011111110101110011110111011011011000101101111110101110101111;
          15:
            level_vec_out = 64'b0100011111110101110011110111011011011000101101111110101110101111;
          16:
            level_vec_out = 64'b0100011111110101110011110111011011011000101101111110101111101111;
          17:
            level_vec_out = 64'b0100011111110111110011110111011011011000101101111110101111101111;
          18:
            level_vec_out = 64'b0100011111110111110111110111011011011000101101111110101111101111;
          19:
            level_vec_out = 64'b0100011111110111110111110111011011011000101111111110101111101111;
          20:
            level_vec_out = 64'b0100011111110111110111111111011111011000101111111111101111111111;
          21:
            level_vec_out = 64'b0100011111110111110111111111011111011000101111111111101111111111;
          22:
            level_vec_out = 64'b0100011111110111110111111111011111011000101111111111101111111111;
          23:
            level_vec_out = 64'b0110011111111111110111111111011111011000101111111111101111111111;
          24:
            level_vec_out = 64'b0110011111111111110111111111011111011000101111111111101111111111;
          25:
            level_vec_out = 64'b0110011111111111110111111111011111011010101111111111101111111111;
          26:
            level_vec_out = 64'b0110011111111111111111111111011111111010111111111111111111111111;
          27:
            level_vec_out = 64'b0110011111111111111111111111011111111011111111111111111111111111;
          28:
            level_vec_out = 64'b0110011111111111111111111111011111111011111111111111111111111111;
          29:
            level_vec_out = 64'b1110011111111111111111111111011111111011111111111111111111111111;
          30:
            level_vec_out = 64'b1110011111111111111111111111011111111111111111111111111111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111011111111111111111111111111111111111;
        endcase
      7:
        case (frame_id)
          0:
            level_vec_out = 64'b0100000110000011111000100000110010001010100000011000111011110101;
          1:
            level_vec_out = 64'b0100000110000011111000100000110010001010100010011000111011110101;
          2:
            level_vec_out = 64'b0100000110000011111000100000110010001010100010011000111011110101;
          3:
            level_vec_out = 64'b0100000110000011111000100000110010001010100010011000111011110101;
          4:
            level_vec_out = 64'b0100000110000011111000100000110010001010100010011000111011110101;
          5:
            level_vec_out = 64'b0100000110000011111001100000110010001010100010011000111011110111;
          6:
            level_vec_out = 64'b0100000110000011111001101000111010001010100011011000111011110111;
          7:
            level_vec_out = 64'b0100000110000011111001101000111010001010100011011000111011110111;
          8:
            level_vec_out = 64'b0100000110010011111001101000111010001010100011011000111011110111;
          9:
            level_vec_out = 64'b0100000110010011111001101000111010001010100111011000111011111111;
          10:
            level_vec_out = 64'b0100000110010011111001101000111010001010100111011000111011111111;
          11:
            level_vec_out = 64'b0101000110010011111001101000111010001010100111011000111111111111;
          12:
            level_vec_out = 64'b0101000110010011111001101000111010101010100111011000111111111111;
          13:
            level_vec_out = 64'b0101000110010011111101101000111010101010100111111000111111111111;
          14:
            level_vec_out = 64'b0101000110010011111101101000111010101110100111111000111111111111;
          15:
            level_vec_out = 64'b1101000110010011111101111000111010101110100111111000111111111111;
          16:
            level_vec_out = 64'b1101000110010011111101111000111010101111100111111000111111111111;
          17:
            level_vec_out = 64'b1101000110010011111101111000111010111111100111111000111111111111;
          18:
            level_vec_out = 64'b1101000110010011111101111000111010111111110111111100111111111111;
          19:
            level_vec_out = 64'b1101000110010111111101111010111010111111110111111100111111111111;
          20:
            level_vec_out = 64'b1101000110011111111101111010111010111111110111111100111111111111;
          21:
            level_vec_out = 64'b1101000111011111111101111010111010111111111111111101111111111111;
          22:
            level_vec_out = 64'b1101000111011111111101111010111110111111111111111101111111111111;
          23:
            level_vec_out = 64'b1101010111011111111101111010111110111111111111111101111111111111;
          24:
            level_vec_out = 64'b1101010111011111111101111010111110111111111111111101111111111111;
          25:
            level_vec_out = 64'b1101010111011111111101111010111110111111111111111101111111111111;
          26:
            level_vec_out = 64'b1101010111011111111101111010111110111111111111111101111111111111;
          27:
            level_vec_out = 64'b1101010111011111111101111010111110111111111111111111111111111111;
          28:
            level_vec_out = 64'b1101010111011111111101111010111110111111111111111111111111111111;
          29:
            level_vec_out = 64'b1111110111011111111101111110111110111111111111111111111111111111;
          30:
            level_vec_out = 64'b1111110111011111111111111110111110111111111111111111111111111111;
          31:
            level_vec_out = 64'b1111110111011111111111111111111111111111111111111111111111111111;
        endcase
    endcase
  end
endmodule