----
 -- @file level_hvec_gen_hdl.hpp
 -- @brief This script generates HDL code for generating high-dimensional LEVEL vectors.
 -- It is a novel method; for more information, please refer to our paper.
 --
 -- @author Saeid Jamili and Marco Angioli
 -- @note Author names are listed in alphabetical order.
 -- @email <saeid.jamili@uniroma1.it>
 -- @email <marco.angioli@uniroma1.it>
 --
 -- @contributors
 --
 -- @date Created: 24th July 2023
 -- @date Last Updated: 23th August 2023
 --
 -- @version 1.0.0
 --
 -- @institute Sapienza University of Rome
 -- @cite https://doi.org/10.xxxx/yyyyy
 --
 -- @section DEPENDENCIES
 -- - Dependency1: Description or version details.
 -- - Dependency2: Description or version details.
 --
 -- @section LICENSE
 -- This file is part of the Aeneas HyperCompute Platform.
 --
 -- Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 --
 -- @section CHANGELOG
 -- @version 1.0.0-dev - 23th August 2023
 -- - Initial release
 --
 -- @todo
 -- - Complete level vector generator function
 -- - Add training
 --
 -- @see
 -- -
 -- -
 -- -
 --
 --

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity level_vec_gen is
    Port ( level_vec_out : out  STD_LOGIC_VECTOR (63 downto 0);
           frame_index : in  STD_LOGIC_VECTOR (2 downto 0);
           frame_id : in  STD_LOGIC_VECTOR (4 downto 0));
end level_vec_gen;

architecture Behavioral of level_vec_gen is
begin
    process (frame_index, frame_id)
    begin
        -- Update this function to match your requirements
        case frame_index is
            when "000" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1110101001000111011010001101101011111000010001010010011000100100";
                    when "00001" => level_vec_out <= "1110101001000111011010001101101011111000010001010010011000100100";
                    when "00010" => level_vec_out <= "1110101001000111011010001101101011111000010001010010011000100100";
                    when "00011" => level_vec_out <= "1110101001000111011010001101101011111010010001010010011000100100";
                    when "00100" => level_vec_out <= "1110101001010111011010101101101011111010010001010010011000101100";
                    when "00101" => level_vec_out <= "1110101001010111011010101101101011111010010001010010011000101110";
                    when "00110" => level_vec_out <= "1110101001011111011010101101101011111010010001011010011000101110";
                    when "00111" => level_vec_out <= "1110101001011111011010101101101011111010010001011010011000101110";
                    when "01000" => level_vec_out <= "1110101001011111011010101101101011111010010001011010011000101110";
                    when "01001" => level_vec_out <= "1110101001011111011010101101101011111110010001011010111000101110";
                    when "01010" => level_vec_out <= "1110101101011111011010111101101011111111010001011110111000101110";
                    when "01011" => level_vec_out <= "1110101101011111011010111101101011111111010001011110111000101110";
                    when "01100" => level_vec_out <= "1110101101011111011010111111101011111111010001011110111000101110";
                    when "01101" => level_vec_out <= "1111101101011111011010111111101011111111010001011110111000101110";
                    when "01110" => level_vec_out <= "1111101101011111111010111111101011111111110001011111111000101110";
                    when "01111" => level_vec_out <= "1111101101011111111010111111101011111111110001011111111000101110";
                    when "10000" => level_vec_out <= "1111101101011111111010111111111011111111111001011111111000101110";
                    when "10001" => level_vec_out <= "1111101101011111111010111111111011111111111001011111111001101110";
                    when "10010" => level_vec_out <= "1111101101011111111010111111111011111111111001011111111001101110";
                    when "10011" => level_vec_out <= "1111101101011111111010111111111011111111111001011111111001101110";
                    when "10100" => level_vec_out <= "1111101101011111111010111111111111111111111001011111111001101110";
                    when "10101" => level_vec_out <= "1111101101011111111010111111111111111111111001111111111001101110";
                    when "10110" => level_vec_out <= "1111101101011111111010111111111111111111111001111111111001101110";
                    when "10111" => level_vec_out <= "1111101101011111111110111111111111111111111001111111111001101110";
                    when "11000" => level_vec_out <= "1111101101011111111110111111111111111111111001111111111001101110";
                    when "11001" => level_vec_out <= "1111101111011111111110111111111111111111111001111111111001101110";
                    when "11010" => level_vec_out <= "1111101111011111111110111111111111111111111101111111111001101110";
                    when "11011" => level_vec_out <= "1111101111011111111110111111111111111111111101111111111101101110";
                    when "11100" => level_vec_out <= "1111101111011111111111111111111111111111111101111111111101101110";
                    when "11101" => level_vec_out <= "1111101111011111111111111111111111111111111101111111111101111110";
                    when "11110" => level_vec_out <= "1111111111011111111111111111111111111111111101111111111101111111";
                    when "11111" => level_vec_out <= "1111111111011111111111111111111111111111111111111111111101111111";
                when others => null;
                end case;
            when "001" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0010100001011000000101101000010011110110100011000100111110100010";
                    when "00001" => level_vec_out <= "0010100001011000000101101000010011110110100011000100111110100010";
                    when "00010" => level_vec_out <= "0010111001111000000101101000010011110110100011000100111110100010";
                    when "00011" => level_vec_out <= "0010111101111000000101101000010011110110100011000100111110100010";
                    when "00100" => level_vec_out <= "0010111101111000000101101000010011110110100011000100111110100010";
                    when "00101" => level_vec_out <= "0011111101111000000101101000010011110110110011000100111110100110";
                    when "00110" => level_vec_out <= "0011111101111000000101101000010011110110110111010110111110100110";
                    when "00111" => level_vec_out <= "0011111101111000000101101000110111110110110111010110111110100110";
                    when "01000" => level_vec_out <= "0011111101111000000101101000110111110110110111010110111110100110";
                    when "01001" => level_vec_out <= "0011111101111000000101101100110111110110110111010110111110100110";
                    when "01010" => level_vec_out <= "0011111101111000000101101100110111110110110111010110111110100110";
                    when "01011" => level_vec_out <= "1011111101111000001101101100110111110110110111010110111110100110";
                    when "01100" => level_vec_out <= "1011111101111000001101101100110111110110110111110110111110110110";
                    when "01101" => level_vec_out <= "1011111101111000001101101100110111110110110111110110111110110110";
                    when "01110" => level_vec_out <= "1011111101111010001101101100110111110110110111110110111110110110";
                    when "01111" => level_vec_out <= "1011111101111010011101101100110111110110110111110110111110110111";
                    when "10000" => level_vec_out <= "1011111101111010011101101110110111110110110111110110111111110111";
                    when "10001" => level_vec_out <= "1011111111111010011101101110110111110110110111110110111111110111";
                    when "10010" => level_vec_out <= "1011111111111010011101101110110111110110111111110111111111110111";
                    when "10011" => level_vec_out <= "1011111111111010011111101110110111110110111111110111111111110111";
                    when "10100" => level_vec_out <= "1011111111111010011111101110110111111110111111110111111111110111";
                    when "10101" => level_vec_out <= "1011111111111010011111101110111111111110111111110111111111110111";
                    when "10110" => level_vec_out <= "1011111111111010111111101110111111111110111111110111111111110111";
                    when "10111" => level_vec_out <= "1011111111111010111111101110111111111110111111110111111111110111";
                    when "11000" => level_vec_out <= "1011111111111011111111101110111111111110111111110111111111110111";
                    when "11001" => level_vec_out <= "1011111111111011111111101110111111111110111111110111111111110111";
                    when "11010" => level_vec_out <= "1011111111111011111111101110111111111110111111110111111111110111";
                    when "11011" => level_vec_out <= "1011111111111011111111101111111111111110111111111111111111110111";
                    when "11100" => level_vec_out <= "1011111111111111111111101111111111111110111111111111111111110111";
                    when "11101" => level_vec_out <= "1011111111111111111111101111111111111110111111111111111111111111";
                    when "11110" => level_vec_out <= "1011111111111111111111101111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111101111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "010" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1101100111011100001000001001010000010101100010010111001000010111";
                    when "00001" => level_vec_out <= "1101100111011100001000001001010000010101100010010111001000010111";
                    when "00010" => level_vec_out <= "1101100111011100001000001001010000010101100010010111001000010111";
                    when "00011" => level_vec_out <= "1101100111011100001000001001010001011101100010010111001000010111";
                    when "00100" => level_vec_out <= "1101100111011100001000001001010001011101100010010111001000110111";
                    when "00101" => level_vec_out <= "1101100111011100001000001001010001011101100010010111011000110111";
                    when "00110" => level_vec_out <= "1101100111011100001010001001010001011101100010010111011000110111";
                    when "00111" => level_vec_out <= "1101100111011101001010001001010001011101100010010111011000110111";
                    when "01000" => level_vec_out <= "1101100111011101001010001101010001011111100010010111011000110111";
                    when "01001" => level_vec_out <= "1101100111011101101010001101010001011111100010010111011000110111";
                    when "01010" => level_vec_out <= "1101100111011101101010001101010001011111100010010111011000110111";
                    when "01011" => level_vec_out <= "1101100111011101101010001101010001011111100010010111011000110111";
                    when "01100" => level_vec_out <= "1101100111011101101010001101010001011111100010010111011001110111";
                    when "01101" => level_vec_out <= "1101100111011101101010001101010001011111100010010111011001110111";
                    when "01110" => level_vec_out <= "1101100111011101101010001101011001011111100010110111011001110111";
                    when "01111" => level_vec_out <= "1101100111011101101010001101011001011111100010110111011001110111";
                    when "10000" => level_vec_out <= "1101100111011101101010001101011001111111100010111111011001110111";
                    when "10001" => level_vec_out <= "1101100111011101101010001101011101111111100010111111011001110111";
                    when "10010" => level_vec_out <= "1101100111011111101010001101011101111111100010111111011001110111";
                    when "10011" => level_vec_out <= "1101100111011111101010001101011101111111100010111111011001110111";
                    when "10100" => level_vec_out <= "1101100111011111101010001101011101111111100010111111011101110111";
                    when "10101" => level_vec_out <= "1101101111011111101010001101011101111111100010111111011101110111";
                    when "10110" => level_vec_out <= "1101101111011111111010001101011111111111100011111111111101110111";
                    when "10111" => level_vec_out <= "1101101111111111111010001101011111111111100011111111111101110111";
                    when "11000" => level_vec_out <= "1101101111111111111011001101011111111111110011111111111111110111";
                    when "11001" => level_vec_out <= "1101101111111111111011001101011111111111110011111111111111111111";
                    when "11010" => level_vec_out <= "1101101111111111111011001101011111111111111011111111111111111111";
                    when "11011" => level_vec_out <= "1111101111111111111011001101011111111111111011111111111111111111";
                    when "11100" => level_vec_out <= "1111101111111111111011001111011111111111111011111111111111111111";
                    when "11101" => level_vec_out <= "1111101111111111111011001111111111111111111111111111111111111111";
                    when "11110" => level_vec_out <= "1111101111111111111111101111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111101111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "011" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1011000101111000101000111010111011110101001000011110011111011111";
                    when "00001" => level_vec_out <= "1011000101111000101000111110111011110101001000011110011111011111";
                    when "00010" => level_vec_out <= "1011000101111000101000111110111011110101001000011110011111011111";
                    when "00011" => level_vec_out <= "1011000101111000101000111110111011110101001000011110011111011111";
                    when "00100" => level_vec_out <= "1011001101111000111000111110111011110101001000011110011111011111";
                    when "00101" => level_vec_out <= "1011001101111000111000111110111011110101001000011110011111011111";
                    when "00110" => level_vec_out <= "1011001101111000111000111110111011110101001000011110011111011111";
                    when "00111" => level_vec_out <= "1011001101111000111000111110111011110101001000011110011111011111";
                    when "01000" => level_vec_out <= "1011101101111000111000111110111011110101001000011111011111011111";
                    when "01001" => level_vec_out <= "1011101101111100111000111110111011110101001000011111011111011111";
                    when "01010" => level_vec_out <= "1011101101111100111000111110111011110101001000011111011111011111";
                    when "01011" => level_vec_out <= "1011101101111100111000111110111011110101001010011111011111011111";
                    when "01100" => level_vec_out <= "1011111101111100111000111110111011110101001010011111011111011111";
                    when "01101" => level_vec_out <= "1111111101111101111000111110111011110101001010011111011111011111";
                    when "01110" => level_vec_out <= "1111111101111101111000111110111011110101001110011111011111011111";
                    when "01111" => level_vec_out <= "1111111101111101111000111110111011110101001110111111011111011111";
                    when "10000" => level_vec_out <= "1111111101111101111010111110111011110101001110111111011111011111";
                    when "10001" => level_vec_out <= "1111111101111101111010111110111011110101101110111111011111111111";
                    when "10010" => level_vec_out <= "1111111101111101111010111110111011110101101110111111111111111111";
                    when "10011" => level_vec_out <= "1111111101111101111010111110111011110111101110111111111111111111";
                    when "10100" => level_vec_out <= "1111111101111101111010111110111011110111101110111111111111111111";
                    when "10101" => level_vec_out <= "1111111101111101111010111110111011110111101111111111111111111111";
                    when "10110" => level_vec_out <= "1111111101111111111010111110111011110111101111111111111111111111";
                    when "10111" => level_vec_out <= "1111111101111111111010111110111011110111101111111111111111111111";
                    when "11000" => level_vec_out <= "1111111101111111111010111110111011111111111111111111111111111111";
                    when "11001" => level_vec_out <= "1111111101111111111010111110111011111111111111111111111111111111";
                    when "11010" => level_vec_out <= "1111111101111111111110111110111111111111111111111111111111111111";
                    when "11011" => level_vec_out <= "1111111101111111111110111110111111111111111111111111111111111111";
                    when "11100" => level_vec_out <= "1111111111111111111110111110111111111111111111111111111111111111";
                    when "11101" => level_vec_out <= "1111111111111111111110111110111111111111111111111111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111110111110111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111110111111111111111111111111111111111111";
                when others => null;
                end case;
            when "100" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1100011101010000111000011110001111010010000101001010110110111000";
                    when "00001" => level_vec_out <= "1100011101010000111000011110001111010010000101001010110110111101";
                    when "00010" => level_vec_out <= "1100011101010000111000011110011111010010000101001010110110111101";
                    when "00011" => level_vec_out <= "1100011101010000111000011110011111010010000101001010110110111101";
                    when "00100" => level_vec_out <= "1100011101010000111000011111011111010010000101001010110110111101";
                    when "00101" => level_vec_out <= "1100011101010000111000011111011111010010000101001010110110111101";
                    when "00110" => level_vec_out <= "1100011101010000111000011111011111010010000101001010110110111101";
                    when "00111" => level_vec_out <= "1100011101010000111000011111011111010010000101101010110111111101";
                    when "01000" => level_vec_out <= "1100011101010000111000011111011111010010000101101010110111111101";
                    when "01001" => level_vec_out <= "1100011101010000111000011111011111010010000101101010110111111101";
                    when "01010" => level_vec_out <= "1100011101010000111000111111011111010010000101101010110111111101";
                    when "01011" => level_vec_out <= "1100011101011000111000111111011111010010000101101110111111111101";
                    when "01100" => level_vec_out <= "1110011101011000111000111111011111010010000101101110111111111101";
                    when "01101" => level_vec_out <= "1110011101011000111000111111011111110010000101101110111111111101";
                    when "01110" => level_vec_out <= "1110011101011000111000111111011111110010000101101110111111111101";
                    when "01111" => level_vec_out <= "1110011101011000111000111111011111110010000101101110111111111101";
                    when "10000" => level_vec_out <= "1110011101011000111000111111011111110010000101101110111111111101";
                    when "10001" => level_vec_out <= "1110011101011000111000111111011111110010000101101110111111111101";
                    when "10010" => level_vec_out <= "1110011101011000111000111111011111110010000101111110111111111101";
                    when "10011" => level_vec_out <= "1110011101111000111000111111111111110010000101111110111111111111";
                    when "10100" => level_vec_out <= "1110011101111000111010111111111111110010010101111110111111111111";
                    when "10101" => level_vec_out <= "1110011101111000111010111111111111110010010101111110111111111111";
                    when "10110" => level_vec_out <= "1110111101111010111010111111111111110010010101111110111111111111";
                    when "10111" => level_vec_out <= "1110111101111010111010111111111111110011010111111110111111111111";
                    when "11000" => level_vec_out <= "1110111101111010111010111111111111110011010111111110111111111111";
                    when "11001" => level_vec_out <= "1110111111111011111010111111111111110011010111111110111111111111";
                    when "11010" => level_vec_out <= "1110111111111011111110111111111111110011010111111110111111111111";
                    when "11011" => level_vec_out <= "1110111111111011111110111111111111110111010111111110111111111111";
                    when "11100" => level_vec_out <= "1111111111111011111110111111111111110111010111111110111111111111";
                    when "11101" => level_vec_out <= "1111111111111011111110111111111111110111010111111111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111110111111111111110111011111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111110111111111111110111111111111111111111111111";
                when others => null;
                end case;
            when "101" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1101110001101000001100011110000101110101101011010001011101001001";
                    when "00001" => level_vec_out <= "1101110001101000001100011110000101110101101011010001011101001011";
                    when "00010" => level_vec_out <= "1101110001101000001100011110000101110101101011010001011101001011";
                    when "00011" => level_vec_out <= "1101110001101000001100011110000101110101101011010001011101001011";
                    when "00100" => level_vec_out <= "1101110001101000001100011110000101110101101011010001011101001011";
                    when "00101" => level_vec_out <= "1101110001101000011100011110000101110101101011010001011101011011";
                    when "00110" => level_vec_out <= "1101110001101000011100011110000101110101101011010001011101011011";
                    when "00111" => level_vec_out <= "1101110001101000011100011110010101110101101011010001011101011011";
                    when "01000" => level_vec_out <= "1101110001101100011100011110010101110101101011010001011101011011";
                    when "01001" => level_vec_out <= "1101110001101100011100011110010101110111101011010001011101011011";
                    when "01010" => level_vec_out <= "1111110001101100011101011110110101110111101011010001011101011011";
                    when "01011" => level_vec_out <= "1111110001101100011101011110110101110111101011010001011101011011";
                    when "01100" => level_vec_out <= "1111110001101100011101011110110101110111101011010001011101011111";
                    when "01101" => level_vec_out <= "1111110001101100011101011110111101110111101011010001011101011111";
                    when "01110" => level_vec_out <= "1111110001101100011101011110111101110111101011010001011101011111";
                    when "01111" => level_vec_out <= "1111110001101100011101011110111101110111101011011001011101011111";
                    when "10000" => level_vec_out <= "1111110001101100011101011110111101110111101011011001011101011111";
                    when "10001" => level_vec_out <= "1111111001101101011101011110111101110111101011011101011101011111";
                    when "10010" => level_vec_out <= "1111111001111101011101011110111101110111101011011111011101011111";
                    when "10011" => level_vec_out <= "1111111001111101011101011110111101110111101011011111111101011111";
                    when "10100" => level_vec_out <= "1111111001111101011101011111111101111111101011011111111101011111";
                    when "10101" => level_vec_out <= "1111111001111101011101011111111101111111101011011111111111011111";
                    when "10110" => level_vec_out <= "1111111001111101011101011111111101111111101011011111111111011111";
                    when "10111" => level_vec_out <= "1111111001111101011101011111111101111111111011011111111111011111";
                    when "11000" => level_vec_out <= "1111111001111101011101011111111101111111111011011111111111011111";
                    when "11001" => level_vec_out <= "1111111001111111011101011111111101111111111111011111111111011111";
                    when "11010" => level_vec_out <= "1111111101111111011101011111111111111111111111011111111111011111";
                    when "11011" => level_vec_out <= "1111111101111111111101011111111111111111111111011111111111011111";
                    when "11100" => level_vec_out <= "1111111101111111111101011111111111111111111111011111111111111111";
                    when "11101" => level_vec_out <= "1111111111111111111101011111111111111111111111011111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111011111111111111111111111011111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111011111111111111111";
                when others => null;
                end case;
            when "110" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1111111101100011010101000001110110010001010011100100000110101001";
                    when "00001" => level_vec_out <= "1111111101100011110101000001110110010011010011100100010110101001";
                    when "00010" => level_vec_out <= "1111111101100011110101000011110110010011010011100100010110101001";
                    when "00011" => level_vec_out <= "1111111101100011110101010011110110010011111011100100010110101001";
                    when "00100" => level_vec_out <= "1111111101100011110101010011110110010011111011100100010110101001";
                    when "00101" => level_vec_out <= "1111111101100011110101010011110110010011111011100100010110101001";
                    when "00110" => level_vec_out <= "1111111101100011110101010111110110010011111011100100010110101001";
                    when "00111" => level_vec_out <= "1111111101100011110101010111110110010011111011100100010110101101";
                    when "01000" => level_vec_out <= "1111111101100011111101010111111110010011111011100100010110101101";
                    when "01001" => level_vec_out <= "1111111101100011111101010111111110011011111011110100010110101101";
                    when "01010" => level_vec_out <= "1111111101100011111101010111111110011011111011110100010110101101";
                    when "01011" => level_vec_out <= "1111111101100011111101010111111110111011111011110100010110111101";
                    when "01100" => level_vec_out <= "1111111101100011111101010111111110111011111011110100010110111101";
                    when "01101" => level_vec_out <= "1111111101100111111101110111111110111011111011110100010110111101";
                    when "01110" => level_vec_out <= "1111111101101111111101110111111110111011111011110100010110111101";
                    when "01111" => level_vec_out <= "1111111101101111111101110111111110111011111011110100010110111101";
                    when "10000" => level_vec_out <= "1111111101101111111101111111111110111011111011110100010110111101";
                    when "10001" => level_vec_out <= "1111111101101111111101111111111110111011111011110100010110111101";
                    when "10010" => level_vec_out <= "1111111101101111111101111111111110111011111011110110010110111101";
                    when "10011" => level_vec_out <= "1111111101101111111101111111111110111011111011110111010110111101";
                    when "10100" => level_vec_out <= "1111111101101111111101111111111110111011111011110111010110111101";
                    when "10101" => level_vec_out <= "1111111101101111111111111111111110111011111011110111110111111101";
                    when "10110" => level_vec_out <= "1111111101101111111111111111111110111011111011110111110111111101";
                    when "10111" => level_vec_out <= "1111111101101111111111111111111110111111111011110111110111111101";
                    when "11000" => level_vec_out <= "1111111101101111111111111111111110111111111011110111110111111101";
                    when "11001" => level_vec_out <= "1111111111101111111111111111111110111111111011110111110111111101";
                    when "11010" => level_vec_out <= "1111111111101111111111111111111111111111111011110111110111111101";
                    when "11011" => level_vec_out <= "1111111111101111111111111111111111111111111011110111110111111111";
                    when "11100" => level_vec_out <= "1111111111111111111111111111111111111111111011110111110111111111";
                    when "11101" => level_vec_out <= "1111111111111111111111111111111111111111111011111111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111111011111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "111" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0100001111011001111011111100100000111101101101111010101101010011";
                    when "00001" => level_vec_out <= "0100001111011001111011111100101000111101101101111010101101010011";
                    when "00010" => level_vec_out <= "0100011111011001111011111100101000111111111101111010101101010011";
                    when "00011" => level_vec_out <= "0100011111011001111011111100101000111111111101111010101111010011";
                    when "00100" => level_vec_out <= "0100011111111001111011111100101000111111111101111010101111010011";
                    when "00101" => level_vec_out <= "0100011111111001111011111100101000111111111101111110101111010011";
                    when "00110" => level_vec_out <= "0100011111111001111011111100111000111111111101111110101111010011";
                    when "00111" => level_vec_out <= "0100011111111001111011111100111001111111111101111110101111010011";
                    when "01000" => level_vec_out <= "0100111111111001111011111100111001111111111101111110101111010011";
                    when "01001" => level_vec_out <= "0100111111111001111011111100111001111111111101111110101111010011";
                    when "01010" => level_vec_out <= "0100111111111001111011111100111001111111111101111110101111010011";
                    when "01011" => level_vec_out <= "0100111111111001111011111100111001111111111101111110101111010011";
                    when "01100" => level_vec_out <= "0100111111111001111111111100111001111111111101111110101111010011";
                    when "01101" => level_vec_out <= "0100111111111011111111111100111001111111111101111110101111010011";
                    when "01110" => level_vec_out <= "0100111111111011111111111100111001111111111101111110101111010011";
                    when "01111" => level_vec_out <= "1100111111111011111111111110111001111111111101111110111111011011";
                    when "10000" => level_vec_out <= "1100111111111011111111111110111001111111111101111110111111011011";
                    when "10001" => level_vec_out <= "1100111111111011111111111110111001111111111101111110111111011011";
                    when "10010" => level_vec_out <= "1100111111111011111111111110111001111111111101111110111111011011";
                    when "10011" => level_vec_out <= "1110111111111011111111111110111001111111111101111110111111011011";
                    when "10100" => level_vec_out <= "1110111111111111111111111110111001111111111101111110111111011011";
                    when "10101" => level_vec_out <= "1110111111111111111111111110111001111111111101111110111111011011";
                    when "10110" => level_vec_out <= "1110111111111111111111111110111001111111111101111110111111011011";
                    when "10111" => level_vec_out <= "1110111111111111111111111110111101111111111101111110111111011111";
                    when "11000" => level_vec_out <= "1110111111111111111111111111111111111111111101111110111111011111";
                    when "11001" => level_vec_out <= "1111111111111111111111111111111111111111111101111110111111011111";
                    when "11010" => level_vec_out <= "1111111111111111111111111111111111111111111101111110111111011111";
                    when "11011" => level_vec_out <= "1111111111111111111111111111111111111111111101111110111111111111";
                    when "11100" => level_vec_out <= "1111111111111111111111111111111111111111111111111110111111111111";
                    when "11101" => level_vec_out <= "1111111111111111111111111111111111111111111111111110111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111111111111110111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when others => null;
        end case;
    end process;
end Behavioral;