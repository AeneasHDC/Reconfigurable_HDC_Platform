----
 -- @file level_hvec_gen_hdl.hpp
 -- @brief This script generates HDL code for generating high-dimensional LEVEL vectors.
 -- It is a novel method; for more information, please refer to our paper.
 --
 -- @author Saeid Jamili and Marco Angioli
 -- @note Author names are listed in alphabetical order.
 -- @email <saeid.jamili@uniroma1.it>
 -- @email <marco.angioli@uniroma1.it>
 --
 -- @contributors
 --
 -- @date Created: 24th July 2023
 -- @date Last Updated: 23th August 2023
 --
 -- @version 1.0.0
 --
 -- @institute Sapienza University of Rome
 -- @cite https://doi.org/10.xxxx/yyyyy
 --
 -- @section DEPENDENCIES
 -- - Dependency1: Description or version details.
 -- - Dependency2: Description or version details.
 --
 -- @section LICENSE
 -- This file is part of the Aeneas HyperCompute Platform.
 --
 -- Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 --
 -- @section CHANGELOG
 -- @version 1.0.0-dev - 23th August 2023
 -- - Initial release
 --
 -- @todo
 -- - Complete level vector generator function
 -- - Add training
 --
 -- @see
 -- -
 -- -
 -- -
 --
 --

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity level_vec_gen is
    Port ( level_vec_out : out  STD_LOGIC_VECTOR (63 downto 0);
           frame_index : in  STD_LOGIC_VECTOR (2 downto 0);
           frame_id : in  STD_LOGIC_VECTOR (4 downto 0));
end level_vec_gen;

architecture Behavioral of level_vec_gen is
begin
    process (frame_index, frame_id)
    begin
        -- Update this function to match your requirements
        case frame_index is
            when "000" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0010010110001110001011101111110000101111010011101100010110001010";
                    when "00001" => level_vec_out <= "0010010110001110001011101111110000101111010011101100010110001010";
                    when "00010" => level_vec_out <= "0010110110001110001011101111110000101111010011101100010110001010";
                    when "00011" => level_vec_out <= "0010110111001110001011101111110000101111010011101100010110001010";
                    when "00100" => level_vec_out <= "0010110111001110001011101111110000101111010011101100010110001010";
                    when "00101" => level_vec_out <= "0010110111001110001011101111110000111111010011101100010110001010";
                    when "00110" => level_vec_out <= "1110110111001110001011101111110000111111011011101100010110001010";
                    when "00111" => level_vec_out <= "1110110111001110001011101111110000111111011011101100010110001010";
                    when "01000" => level_vec_out <= "1110110111001110001011101111111000111111011011101100010110001110";
                    when "01001" => level_vec_out <= "1110110111001110001011101111111000111111011011101100010111001110";
                    when "01010" => level_vec_out <= "1110110111001110001011101111111000111111011011101100110111001110";
                    when "01011" => level_vec_out <= "1110110111001110001011101111111000111111011011101100110111001111";
                    when "01100" => level_vec_out <= "1110110111001110001011111111111000111111011011101100110111001111";
                    when "01101" => level_vec_out <= "1110110111001110001011111111111000111111011011101110110111001111";
                    when "01110" => level_vec_out <= "1110110111001110001011111111111000111111011011101110110111011111";
                    when "01111" => level_vec_out <= "1110110111001110101011111111111000111111011011101110110111011111";
                    when "10000" => level_vec_out <= "1110110111101110101011111111111000111111011011101110110111111111";
                    when "10001" => level_vec_out <= "1110110111101110101011111111111010111111011111101110110111111111";
                    when "10010" => level_vec_out <= "1110110111101110101011111111111010111111011111111110111111111111";
                    when "10011" => level_vec_out <= "1110110111101110101011111111111010111111011111111110111111111111";
                    when "10100" => level_vec_out <= "1110110111101110101011111111111010111111011111111110111111111111";
                    when "10101" => level_vec_out <= "1110110111101110101011111111111010111111011111111110111111111111";
                    when "10110" => level_vec_out <= "1110110111101110101011111111111010111111111111111111111111111111";
                    when "10111" => level_vec_out <= "1110110111101111101011111111111010111111111111111111111111111111";
                    when "11000" => level_vec_out <= "1110110111101111101011111111111011111111111111111111111111111111";
                    when "11001" => level_vec_out <= "1110110111101111101011111111111011111111111111111111111111111111";
                    when "11010" => level_vec_out <= "1110111111111111101011111111111011111111111111111111111111111111";
                    when "11011" => level_vec_out <= "1110111111111111101011111111111011111111111111111111111111111111";
                    when "11100" => level_vec_out <= "1110111111111111101111111111111011111111111111111111111111111111";
                    when "11101" => level_vec_out <= "1111111111111111101111111111111011111111111111111111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111101111111111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111101111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "001" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0011100000010100100000100011100100011110001101110001111111111100";
                    when "00001" => level_vec_out <= "0011100000010100100000100011100100011110001101110001111111111101";
                    when "00010" => level_vec_out <= "0011100000010100100010100011100100011110011101110001111111111101";
                    when "00011" => level_vec_out <= "0011100001010100100010100011100100011110011101110001111111111101";
                    when "00100" => level_vec_out <= "0011100001010110100110100011100100011110011101110001111111111101";
                    when "00101" => level_vec_out <= "0011100001110110100110100011100100011110011101110001111111111101";
                    when "00110" => level_vec_out <= "0011100001110110100110100011100100011110011101110001111111111101";
                    when "00111" => level_vec_out <= "0011100001110110100110100011100100011110011101110001111111111101";
                    when "01000" => level_vec_out <= "0011100001110110100110100011100100011110011101110001111111111101";
                    when "01001" => level_vec_out <= "0011100001110110100110100011110100011110011111110001111111111101";
                    when "01010" => level_vec_out <= "0011100001110110100110101011111100011110011111110001111111111101";
                    when "01011" => level_vec_out <= "0011101001110110100110101011111100011110011111110001111111111101";
                    when "01100" => level_vec_out <= "0011101001110110100110101011111100111110011111110001111111111101";
                    when "01101" => level_vec_out <= "0011101001110110100110101011111100111110011111110001111111111101";
                    when "01110" => level_vec_out <= "0011101001110110100110101011111100111110111111110001111111111101";
                    when "01111" => level_vec_out <= "0011101001110110100110101011111101111110111111110001111111111101";
                    when "10000" => level_vec_out <= "0011101001110110100110101011111101111110111111110001111111111101";
                    when "10001" => level_vec_out <= "0011101001110110100110101111111101111110111111110001111111111101";
                    when "10010" => level_vec_out <= "0011101011111110100110111111111101111110111111110011111111111101";
                    when "10011" => level_vec_out <= "0111101011111110100110111111111101111111111111111011111111111101";
                    when "10100" => level_vec_out <= "0111101011111110100110111111111101111111111111111011111111111101";
                    when "10101" => level_vec_out <= "0111101111111110100110111111111101111111111111111011111111111101";
                    when "10110" => level_vec_out <= "0111101111111110100110111111111101111111111111111011111111111101";
                    when "10111" => level_vec_out <= "0111101111111110100110111111111101111111111111111011111111111101";
                    when "11000" => level_vec_out <= "0111101111111110100110111111111101111111111111111011111111111101";
                    when "11001" => level_vec_out <= "0111101111111110110110111111111101111111111111111011111111111101";
                    when "11010" => level_vec_out <= "1111101111111110110110111111111101111111111111111011111111111101";
                    when "11011" => level_vec_out <= "1111101111111111110110111111111101111111111111111011111111111101";
                    when "11100" => level_vec_out <= "1111101111111111110111111111111111111111111111111011111111111101";
                    when "11101" => level_vec_out <= "1111101111111111110111111111111111111111111111111111111111111101";
                    when "11110" => level_vec_out <= "1111111111111111110111111111111111111111111111111111111111111101";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111101";
                when others => null;
                end case;
            when "010" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1001111111110010110001101100111110110000011010111101010110111110";
                    when "00001" => level_vec_out <= "1001111111110010110001101100111110110000011010111101010110111110";
                    when "00010" => level_vec_out <= "1001111111110010110001101100111110110000011010111101010110111110";
                    when "00011" => level_vec_out <= "1001111111110010110001101100111110110010011010111101010110111110";
                    when "00100" => level_vec_out <= "1001111111110010110001111100111110110010011010111101010110111110";
                    when "00101" => level_vec_out <= "1001111111110010110001111100111110110010011010111101010110111110";
                    when "00110" => level_vec_out <= "1001111111110010110001111100111111110010011010111101010110111110";
                    when "00111" => level_vec_out <= "1001111111110010110001111100111111110010111010111101010110111110";
                    when "01000" => level_vec_out <= "1001111111110010111001111100111111110010111010111101010110111110";
                    when "01001" => level_vec_out <= "1001111111110010111001111110111111110010111010111101010110111110";
                    when "01010" => level_vec_out <= "1001111111110010111001111110111111110010111010111101010110111110";
                    when "01011" => level_vec_out <= "1001111111110010111001111110111111110010111010111111010110111110";
                    when "01100" => level_vec_out <= "1001111111110010111101111110111111110010111010111111010110111110";
                    when "01101" => level_vec_out <= "1001111111110010111101111110111111110010111110111111010110111110";
                    when "01110" => level_vec_out <= "1101111111110010111101111110111111111010111110111111011110111110";
                    when "01111" => level_vec_out <= "1101111111110010111101111110111111111010111110111111011111111111";
                    when "10000" => level_vec_out <= "1101111111110010111101111110111111111010111110111111011111111111";
                    when "10001" => level_vec_out <= "1101111111110010111101111110111111111010111111111111011111111111";
                    when "10010" => level_vec_out <= "1101111111110010111101111110111111111010111111111111011111111111";
                    when "10011" => level_vec_out <= "1101111111110011111101111110111111111010111111111111011111111111";
                    when "10100" => level_vec_out <= "1101111111110011111101111111111111111010111111111111011111111111";
                    when "10101" => level_vec_out <= "1101111111110011111101111111111111111010111111111111011111111111";
                    when "10110" => level_vec_out <= "1101111111110011111101111111111111111010111111111111011111111111";
                    when "10111" => level_vec_out <= "1101111111110111111101111111111111111010111111111111011111111111";
                    when "11000" => level_vec_out <= "1101111111110111111101111111111111111010111111111111011111111111";
                    when "11001" => level_vec_out <= "1101111111110111111101111111111111111110111111111111011111111111";
                    when "11010" => level_vec_out <= "1101111111110111111111111111111111111110111111111111011111111111";
                    when "11011" => level_vec_out <= "1101111111110111111111111111111111111110111111111111011111111111";
                    when "11100" => level_vec_out <= "1101111111110111111111111111111111111110111111111111011111111111";
                    when "11101" => level_vec_out <= "1101111111111111111111111111111111111110111111111111011111111111";
                    when "11110" => level_vec_out <= "1101111111111111111111111111111111111110111111111111011111111111";
                    when "11111" => level_vec_out <= "1101111111111111111111111111111111111111111111111111011111111111";
                when others => null;
                end case;
            when "011" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1001100011001001010000100101101001100011010100100111100110000001";
                    when "00001" => level_vec_out <= "1001100011001001010100100101101001100111010100100111101110001001";
                    when "00010" => level_vec_out <= "1001100011001001110100100101101001100111010100100111101110001001";
                    when "00011" => level_vec_out <= "1001100011001101110100100101101001100111010100100111101110001001";
                    when "00100" => level_vec_out <= "1001100011001101110100100101111001100111010100100111111110001001";
                    when "00101" => level_vec_out <= "1001100011001101110100100101111101100111010101100111111110001001";
                    when "00110" => level_vec_out <= "1001100111001101110100100101111101100111010101100111111110001001";
                    when "00111" => level_vec_out <= "1001100111101101110100100101111101100111010101100111111110001001";
                    when "01000" => level_vec_out <= "1001100111101101110100100101111101100111010101100111111110001001";
                    when "01001" => level_vec_out <= "1001100111101101111100100111111101100111010101100111111110001001";
                    when "01010" => level_vec_out <= "1001100111101101111100100111111101100111010101100111111110001001";
                    when "01011" => level_vec_out <= "1001100111101101111100100111111101100111110101100111111110001001";
                    when "01100" => level_vec_out <= "1101100111101101111100100111111101100111110101100111111110001001";
                    when "01101" => level_vec_out <= "1101100111101101111110100111111101100111110101110111111110101001";
                    when "01110" => level_vec_out <= "1101100111101101111110100111111101100111110101110111111110101001";
                    when "01111" => level_vec_out <= "1101101111101101111110100111111101100111110101110111111110101001";
                    when "10000" => level_vec_out <= "1101101111101101111110100111111101100111110101110111111110101101";
                    when "10001" => level_vec_out <= "1101101111101101111110100111111101100111110101110111111110101101";
                    when "10010" => level_vec_out <= "1101101111101101111110100111111101100111110101110111111110101101";
                    when "10011" => level_vec_out <= "1101101111101101111110110111111101100111110101110111111110101101";
                    when "10100" => level_vec_out <= "1101101111101101111110110111111101100111110101110111111110111101";
                    when "10101" => level_vec_out <= "1101111111101101111110110111111101100111110101110111111110111101";
                    when "10110" => level_vec_out <= "1101111111101101111110110111111101100111110101110111111110111101";
                    when "10111" => level_vec_out <= "1101111111101101111110110111111101100111111101110111111111111101";
                    when "11000" => level_vec_out <= "1101111111101111111110110111111101100111111101111111111111111111";
                    when "11001" => level_vec_out <= "1101111111101111111110111111111101100111111101111111111111111111";
                    when "11010" => level_vec_out <= "1101111111101111111110111111111101100111111101111111111111111111";
                    when "11011" => level_vec_out <= "1101111111101111111110111111111101110111111111111111111111111111";
                    when "11100" => level_vec_out <= "1101111111111111111111111111111101111111111111111111111111111111";
                    when "11101" => level_vec_out <= "1101111111111111111111111111111111111111111111111111111111111111";
                    when "11110" => level_vec_out <= "1101111111111111111111111111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1101111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "100" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0001011110101100001111000100111001110101011111001111101101011011";
                    when "00001" => level_vec_out <= "0001011110101100001111000100111001110101011111001111101101011111";
                    when "00010" => level_vec_out <= "0001011110101100001111000100111011110101011111001111101101011111";
                    when "00011" => level_vec_out <= "0001011110101100001111000100111011110101011111001111101101011111";
                    when "00100" => level_vec_out <= "0001011110101100001111000100111011110111011111001111101101011111";
                    when "00101" => level_vec_out <= "0001011110101101001111000100111011110111111111001111101101011111";
                    when "00110" => level_vec_out <= "0001011110101101001111000110111011110111111111001111101101011111";
                    when "00111" => level_vec_out <= "0001011110101101001111000110111011110111111111001111101101011111";
                    when "01000" => level_vec_out <= "0001011110101101001111000110111011110111111111001111101101011111";
                    when "01001" => level_vec_out <= "0001011110101101001111000110111011110111111111001111101101011111";
                    when "01010" => level_vec_out <= "0001011111101101001111000110111111110111111111001111101101011111";
                    when "01011" => level_vec_out <= "0001011111101101001111000110111111110111111111001111101101011111";
                    when "01100" => level_vec_out <= "0001011111101101001111000110111111110111111111001111101101011111";
                    when "01101" => level_vec_out <= "0001011111101101001111000110111111110111111111001111101101011111";
                    when "01110" => level_vec_out <= "0001011111101101001111000110111111110111111111001111101101011111";
                    when "01111" => level_vec_out <= "0011011111101101001111000110111111110111111111001111101101011111";
                    when "10000" => level_vec_out <= "0011011111101101001111000110111111110111111111001111101101011111";
                    when "10001" => level_vec_out <= "0011011111101101001111100111111111110111111111001111101101011111";
                    when "10010" => level_vec_out <= "0011011111101101001111100111111111110111111111001111101101011111";
                    when "10011" => level_vec_out <= "0011011111101101001111100111111111110111111111001111101101011111";
                    when "10100" => level_vec_out <= "0011011111101101001111100111111111110111111111001111111101011111";
                    when "10101" => level_vec_out <= "0011011111101101001111100111111111110111111111001111111101011111";
                    when "10110" => level_vec_out <= "0011011111101101111111100111111111110111111111001111111101011111";
                    when "10111" => level_vec_out <= "0011011111101101111111100111111111110111111111001111111101111111";
                    when "11000" => level_vec_out <= "0011011111101101111111100111111111110111111111001111111101111111";
                    when "11001" => level_vec_out <= "0011011111101101111111100111111111110111111111101111111101111111";
                    when "11010" => level_vec_out <= "0011011111111101111111110111111111110111111111101111111101111111";
                    when "11011" => level_vec_out <= "1111011111111111111111110111111111110111111111101111111101111111";
                    when "11100" => level_vec_out <= "1111011111111111111111110111111111111111111111101111111101111111";
                    when "11101" => level_vec_out <= "1111011111111111111111110111111111111111111111101111111101111111";
                    when "11110" => level_vec_out <= "1111011111111111111111111111111111111111111111101111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "101" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0101101001100110100110000010011001011111011110110100110101001100";
                    when "00001" => level_vec_out <= "0101101001110110100110000010011001011111011110110100110101001100";
                    when "00010" => level_vec_out <= "0101101001110110100110000010011101011111011110110100110101001100";
                    when "00011" => level_vec_out <= "0101101001110110100110000010011101011111011110110100110101001100";
                    when "00100" => level_vec_out <= "0101101001110110100110000010011101011111011110110100110101001100";
                    when "00101" => level_vec_out <= "0101111001110110100110000010011101011111011110110100110101001100";
                    when "00110" => level_vec_out <= "0101111001110110100110000010011101011111011110110100110101001100";
                    when "00111" => level_vec_out <= "0101111001110110110110001010011101011111011110110100110101001100";
                    when "01000" => level_vec_out <= "0111111001110110110110001011011101011111011110110100110101101100";
                    when "01001" => level_vec_out <= "1111111001110110110110001011011101011111011110110100110101101100";
                    when "01010" => level_vec_out <= "1111111001110110110110011011011101011111011110110100110101101110";
                    when "01011" => level_vec_out <= "1111111001110110110110111011011101011111011110110100110111101110";
                    when "01100" => level_vec_out <= "1111111001110110110110111011011101011111011110110101110111101110";
                    when "01101" => level_vec_out <= "1111111001110110110110111111011101011111011110110101110111101110";
                    when "01110" => level_vec_out <= "1111111001110110110110111111011111011111011110110101110111111110";
                    when "01111" => level_vec_out <= "1111111001110110110110111111011111011111011110110101110111111110";
                    when "10000" => level_vec_out <= "1111111001110110110110111111011111011111011110111101110111111110";
                    when "10001" => level_vec_out <= "1111111001110110110111111111011111011111011110111101110111111110";
                    when "10010" => level_vec_out <= "1111111001110110110111111111011111011111011110111101110111111110";
                    when "10011" => level_vec_out <= "1111111001110110110111111111011111111111011110111111110111111110";
                    when "10100" => level_vec_out <= "1111111101110110110111111111111111111111011110111111110111111110";
                    when "10101" => level_vec_out <= "1111111111110110110111111111111111111111011110111111110111111110";
                    when "10110" => level_vec_out <= "1111111111110110110111111111111111111111011110111111110111111110";
                    when "10111" => level_vec_out <= "1111111111110110110111111111111111111111011110111111110111111110";
                    when "11000" => level_vec_out <= "1111111111110110110111111111111111111111011110111111111111111110";
                    when "11001" => level_vec_out <= "1111111111110110110111111111111111111111011111111111111111111110";
                    when "11010" => level_vec_out <= "1111111111110111110111111111111111111111011111111111111111111110";
                    when "11011" => level_vec_out <= "1111111111111111111111111111111111111111011111111111111111111110";
                    when "11100" => level_vec_out <= "1111111111111111111111111111111111111111011111111111111111111110";
                    when "11101" => level_vec_out <= "1111111111111111111111111111111111111111011111111111111111111110";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111011111111111111111111110";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111011111111111111111111111";
                when others => null;
                end case;
            when "110" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1101010000000111000100110011110000100010111100000100111001101100";
                    when "00001" => level_vec_out <= "1101010000000111000100110011110000100010111100000100111001101100";
                    when "00010" => level_vec_out <= "1101010000000111000100110111110000100110111100000100111001101100";
                    when "00011" => level_vec_out <= "1101010100000111000100110111110000100110111100000100111101101100";
                    when "00100" => level_vec_out <= "1101010100000111000100110111110000100110111100000110111111101100";
                    when "00101" => level_vec_out <= "1101010100000111000100110111110000100110111100000110111111101100";
                    when "00110" => level_vec_out <= "1101010110000111000100110111110000100110111100000110111111101100";
                    when "00111" => level_vec_out <= "1111010110000111000100110111110000100110111100000110111111101100";
                    when "01000" => level_vec_out <= "1111010110000111000100110111110000100110111100000110111111101101";
                    when "01001" => level_vec_out <= "1111010110000111000100110111110000100110111110000110111111101101";
                    when "01010" => level_vec_out <= "1111010110000111000101110111110000100110111110000110111111101101";
                    when "01011" => level_vec_out <= "1111010110000111000101110111110100100110111110000110111111101101";
                    when "01100" => level_vec_out <= "1111010110001111000101110111110101100110111110000110111111101101";
                    when "01101" => level_vec_out <= "1111010110011111000101110111110101101110111110000110111111101101";
                    when "01110" => level_vec_out <= "1111010110011111000101110111110101101110111110000110111111101101";
                    when "01111" => level_vec_out <= "1111010110011111000101110111110101101110111110001110111111101101";
                    when "10000" => level_vec_out <= "1111010110011111000101110111110101101110111110001110111111101101";
                    when "10001" => level_vec_out <= "1111010110011111000101110111110101101110111111001110111111101101";
                    when "10010" => level_vec_out <= "1111010110011111000101110111111101101110111111001110111111101111";
                    when "10011" => level_vec_out <= "1111010111011111000101110111111101101110111111001110111111101111";
                    when "10100" => level_vec_out <= "1111010111011111000101110111111101101110111111001110111111101111";
                    when "10101" => level_vec_out <= "1111110111011111000101110111111101111110111111001110111111101111";
                    when "10110" => level_vec_out <= "1111110111011111000101111111111111111110111111001110111111101111";
                    when "10111" => level_vec_out <= "1111110111011111100101111111111111111110111111001111111111101111";
                    when "11000" => level_vec_out <= "1111110111011111100111111111111111111110111111001111111111101111";
                    when "11001" => level_vec_out <= "1111110111011111110111111111111111111110111111011111111111101111";
                    when "11010" => level_vec_out <= "1111110111011111111111111111111111111110111111011111111111101111";
                    when "11011" => level_vec_out <= "1111110111011111111111111111111111111110111111011111111111101111";
                    when "11100" => level_vec_out <= "1111111111011111111111111111111111111110111111011111111111101111";
                    when "11101" => level_vec_out <= "1111111111011111111111111111111111111110111111011111111111101111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111111111011111111111101111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111011111111111111111";
                when others => null;
                end case;
            when "111" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1001110100000101000100110110101000010000000110011011100000101101";
                    when "00001" => level_vec_out <= "1001110100000101000100110110101010010000000110011011100000101101";
                    when "00010" => level_vec_out <= "1001110100000101000100110110101010010000000110011011100000101101";
                    when "00011" => level_vec_out <= "1101111100000101000100110110101010010000000110011011100000101101";
                    when "00100" => level_vec_out <= "1101111100000101000100110110101010010000000110011011100000101101";
                    when "00101" => level_vec_out <= "1101111100000101000100110110101010010000000110011111100000101101";
                    when "00110" => level_vec_out <= "1101111100000101000100110110101010010000000110011111100000101111";
                    when "00111" => level_vec_out <= "1101111100000101000100111110101110010000000110011111100001101111";
                    when "01000" => level_vec_out <= "1101111100000101000100111110101110010000100110011111100001101111";
                    when "01001" => level_vec_out <= "1101111100000101000100111110101110010000100110011111100001101111";
                    when "01010" => level_vec_out <= "1101111100000101000100111110101110010000100110011111100001101111";
                    when "01011" => level_vec_out <= "1101111100000101000100111110101110010000100110011111101001101111";
                    when "01100" => level_vec_out <= "1111111100000101000100111110101110010000100110011111101001101111";
                    when "01101" => level_vec_out <= "1111111100000101000100111110101110010000100110011111101001101111";
                    when "01110" => level_vec_out <= "1111111100000101000100111110101110010000100111011111101001101111";
                    when "01111" => level_vec_out <= "1111111100000101000100111110101111010000100111011111101001101111";
                    when "10000" => level_vec_out <= "1111111100010101000100111111101111010010101111011111101001101111";
                    when "10001" => level_vec_out <= "1111111100010101000100111111101111010010101111011111101001101111";
                    when "10010" => level_vec_out <= "1111111100010101000100111111101111010010101111011111101001101111";
                    when "10011" => level_vec_out <= "1111111100010101000100111111101111010010101111011111101001101111";
                    when "10100" => level_vec_out <= "1111111110010101000100111111101111010010101111111111101001111111";
                    when "10101" => level_vec_out <= "1111111110010101010101111111111111010010101111111111101001111111";
                    when "10110" => level_vec_out <= "1111111111010101010101111111111111010011101111111111101001111111";
                    when "10111" => level_vec_out <= "1111111111010101010101111111111111110011101111111111101001111111";
                    when "11000" => level_vec_out <= "1111111111010101011101111111111111111011101111111111101001111111";
                    when "11001" => level_vec_out <= "1111111111010101011101111111111111111011101111111111101011111111";
                    when "11010" => level_vec_out <= "1111111111010101011101111111111111111011101111111111101011111111";
                    when "11011" => level_vec_out <= "1111111111010101011101111111111111111011101111111111101011111111";
                    when "11100" => level_vec_out <= "1111111111010101011101111111111111111011101111111111101011111111";
                    when "11101" => level_vec_out <= "1111111111010101111101111111111111111111111111111111111011111111";
                    when "11110" => level_vec_out <= "1111111111111101111101111111111111111111111111111111111011111111";
                    when "11111" => level_vec_out <= "1111111111111101111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when others => null;
        end case;
    end process;
end Behavioral;