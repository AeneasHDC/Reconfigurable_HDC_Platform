----
 -- @file level_hvec_gen_hdl.hpp
 -- @brief This script generates HDL code for generating high-dimensional LEVEL vectors.
 -- It is a novel method; for more information, please refer to our paper.
 --
 -- @author Saeid Jamili and Marco Angioli
 -- @note Author names are listed in alphabetical order.
 -- @email <saeid.jamili@uniroma1.it>
 -- @email <marco.angioli@uniroma1.it>
 --
 -- @contributors
 --
 -- @date Created: 24th July 2023
 -- @date Last Updated: 23th August 2023
 --
 -- @version 1.0.0
 --
 -- @institute Sapienza University of Rome
 -- @cite https://doi.org/10.xxxx/yyyyy
 --
 -- @section DEPENDENCIES
 -- - Dependency1: Description or version details.
 -- - Dependency2: Description or version details.
 --
 -- @section LICENSE
 -- This file is part of the Aeneas HyperCompute Platform.
 --
 -- Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 --
 -- @section CHANGELOG
 -- @version 1.0.0-dev - 23th August 2023
 -- - Initial release
 --
 -- @todo
 -- - Complete level vector generator function
 -- - Add training
 --
 -- @see
 -- -
 -- -
 -- -
 --
 --

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity level_vec_gen is
    Port ( level_vec_out : out  STD_LOGIC_VECTOR (63 downto 0);
           frame_index : in  STD_LOGIC_VECTOR (2 downto 0);
           frame_id : in  STD_LOGIC_VECTOR (4 downto 0));
end level_vec_gen;

architecture Behavioral of level_vec_gen is
begin
    process (frame_index, frame_id)
    begin
        -- Update this function to match your requirements
        case frame_index is
            when "000" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1100111110100110001101001001101011111110001110010011011001100000";
                    when "00001" => level_vec_out <= "1100111110100110001101001001101011111110001111010011011101100000";
                    when "00010" => level_vec_out <= "1100111110100110011101001001101011111110101111010011011101100000";
                    when "00011" => level_vec_out <= "1100111110100110011101001001101011111110101111010011011101100000";
                    when "00100" => level_vec_out <= "1100111110100110011101001001101011111110101111010111011101100000";
                    when "00101" => level_vec_out <= "1100111110100110011101001001101011111110101111010111011101100000";
                    when "00110" => level_vec_out <= "1100111110100110011101001001101011111110101111010111011101100000";
                    when "00111" => level_vec_out <= "1100111111100110011101001001101011111110101111010111011101100000";
                    when "01000" => level_vec_out <= "1100111111100110011101001001101111111110101111010111011101100000";
                    when "01001" => level_vec_out <= "1100111111100110011101001001101111111110101111010111011101100000";
                    when "01010" => level_vec_out <= "1101111111110110011101001001101111111110101111010111011101100000";
                    when "01011" => level_vec_out <= "1101111111110110011101001001101111111110101111010111011101100000";
                    when "01100" => level_vec_out <= "1101111111110110011101001001101111111110101111010111111101100000";
                    when "01101" => level_vec_out <= "1101111111110110011101001001101111111110101111010111111101100000";
                    when "01110" => level_vec_out <= "1101111111110110111101001001101111111110111111010111111101100000";
                    when "01111" => level_vec_out <= "1101111111110110111101001001101111111110111111010111111101100000";
                    when "10000" => level_vec_out <= "1101111111110110111101001001101111111110111111010111111101110000";
                    when "10001" => level_vec_out <= "1101111111110110111101001001101111111110111111010111111101111000";
                    when "10010" => level_vec_out <= "1101111111110110111101001001101111111110111111110111111101111000";
                    when "10011" => level_vec_out <= "1101111111110110111101001001101111111110111111110111111101111000";
                    when "10100" => level_vec_out <= "1101111111110110111101001001101111111111111111110111111101111001";
                    when "10101" => level_vec_out <= "1101111111110110111101001001101111111111111111110111111101111011";
                    when "10110" => level_vec_out <= "1101111111110110111101001001101111111111111111110111111101111011";
                    when "10111" => level_vec_out <= "1101111111110110111101001001101111111111111111110111111101111011";
                    when "11000" => level_vec_out <= "1101111111110110111101001001101111111111111111110111111101111011";
                    when "11001" => level_vec_out <= "1101111111110110111101001001101111111111111111110111111111111011";
                    when "11010" => level_vec_out <= "1101111111110110111101001001101111111111111111110111111111111111";
                    when "11011" => level_vec_out <= "1101111111110110111101001001111111111111111111110111111111111111";
                    when "11100" => level_vec_out <= "1101111111110110111101001001111111111111111111110111111111111111";
                    when "11101" => level_vec_out <= "1101111111111110111101101011111111111111111111110111111111111111";
                    when "11110" => level_vec_out <= "1101111111111110111101111111111111111111111111110111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111101111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "001" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0100000101100111011001010111101111001001001111010010011100100110";
                    when "00001" => level_vec_out <= "0100000101100111011001010111101111001001001111010010011100100110";
                    when "00010" => level_vec_out <= "0100001111100111011001010111101111001001001111010011011100100110";
                    when "00011" => level_vec_out <= "0100001111100111011001010111111111001001001111010011011100100110";
                    when "00100" => level_vec_out <= "0100001111100111011001011111111111001001001111010011011100100110";
                    when "00101" => level_vec_out <= "0100001111100111011001011111111111011001001111010011011100100110";
                    when "00110" => level_vec_out <= "0100001111100111011001011111111111011001001111010011011100100110";
                    when "00111" => level_vec_out <= "0100001111100111011001011111111111011001001111010011011100100110";
                    when "01000" => level_vec_out <= "0100001111100111011011011111111111011001001111010011011100100110";
                    when "01001" => level_vec_out <= "0100001111100111011011011111111111011001001111010011011100100110";
                    when "01010" => level_vec_out <= "0100001111100111011011011111111111011001001111010011111100100110";
                    when "01011" => level_vec_out <= "0100001111100111011011011111111111011001001111010011111100100110";
                    when "01100" => level_vec_out <= "0100001111100111011111011111111111011001001111110011111101100110";
                    when "01101" => level_vec_out <= "0100001111100111011111011111111111011001001111110011111101100110";
                    when "01110" => level_vec_out <= "0100001111100111011111011111111111011001001111110011111101100110";
                    when "01111" => level_vec_out <= "0110001111100111011111011111111111011001001111110011111101100110";
                    when "10000" => level_vec_out <= "0110001111100111011111011111111111011001001111110011111101100110";
                    when "10001" => level_vec_out <= "0111101111100111011111011111111111011001001111110011111101101110";
                    when "10010" => level_vec_out <= "0111101111100111111111011111111111011001001111110011111101101110";
                    when "10011" => level_vec_out <= "0111101111100111111111011111111111011001001111110011111101101110";
                    when "10100" => level_vec_out <= "0111101111100111111111011111111111011001001111111011111101101110";
                    when "10101" => level_vec_out <= "0111101111110111111111011111111111011001011111111011111101101110";
                    when "10110" => level_vec_out <= "0111101111111111111111011111111111011001011111111011111101101110";
                    when "10111" => level_vec_out <= "0111101111111111111111111111111111111001011111111011111101101111";
                    when "11000" => level_vec_out <= "0111101111111111111111111111111111111001111111111011111101101111";
                    when "11001" => level_vec_out <= "0111101111111111111111111111111111111101111111111011111101101111";
                    when "11010" => level_vec_out <= "0111101111111111111111111111111111111101111111111111111101101111";
                    when "11011" => level_vec_out <= "0111101111111111111111111111111111111111111111111111111101101111";
                    when "11100" => level_vec_out <= "0111101111111111111111111111111111111111111111111111111101111111";
                    when "11101" => level_vec_out <= "0111111111111111111111111111111111111111111111111111111111111111";
                    when "11110" => level_vec_out <= "0111111111111111111111111111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "0111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "010" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0110001011000101101011110000001100110001110111000000010001001011";
                    when "00001" => level_vec_out <= "0110001011000101101011110000001100110001110111000000010001001011";
                    when "00010" => level_vec_out <= "0110001011000101101011110000001100110001110111000000010001001011";
                    when "00011" => level_vec_out <= "0110001011010101101011110000001100110001110111000000010001001011";
                    when "00100" => level_vec_out <= "0110001011010101101011110000001100110001110111000000010001011011";
                    when "00101" => level_vec_out <= "0111001111010101101011110000001100110001110111000000010001011011";
                    when "00110" => level_vec_out <= "0111001111010101101011110100001100110001111111000010010001011011";
                    when "00111" => level_vec_out <= "0111011111010101101011110100001100110001111111000010010001011011";
                    when "01000" => level_vec_out <= "0111111111010101101011110100001100110001111111000010010001011011";
                    when "01001" => level_vec_out <= "0111111111110111101011110100001100110101111111000010010001011011";
                    when "01010" => level_vec_out <= "0111111111110111101011110100001100110101111111000010010001011011";
                    when "01011" => level_vec_out <= "0111111111110111101011110110001100110101111111000010010001011011";
                    when "01100" => level_vec_out <= "0111111111110111101011110110001100110101111111000010010001011011";
                    when "01101" => level_vec_out <= "0111111111110111101011110110011100110101111111000010010001011011";
                    when "01110" => level_vec_out <= "0111111111110111101011110110011100110101111111000010010001011111";
                    when "01111" => level_vec_out <= "1111111111110111101011110110011100110101111111000010010001011111";
                    when "10000" => level_vec_out <= "1111111111110111101011110110011101110101111111000010011001011111";
                    when "10001" => level_vec_out <= "1111111111110111101011110110011101110101111111000010011001011111";
                    when "10010" => level_vec_out <= "1111111111110111101011110110011101110111111111000010011001011111";
                    when "10011" => level_vec_out <= "1111111111110111101011110110011111110111111111000010011001011111";
                    when "10100" => level_vec_out <= "1111111111110111101011110110011111110111111111010110011001011111";
                    when "10101" => level_vec_out <= "1111111111110111101011110110011111111111111111010110011001011111";
                    when "10110" => level_vec_out <= "1111111111111111101011110110011111111111111111010110011001011111";
                    when "10111" => level_vec_out <= "1111111111111111101011110110011111111111111111010110011001111111";
                    when "11000" => level_vec_out <= "1111111111111111101011110110011111111111111111010110111011111111";
                    when "11001" => level_vec_out <= "1111111111111111101011110111011111111111111111011110111011111111";
                    when "11010" => level_vec_out <= "1111111111111111101011110111011111111111111111011110111011111111";
                    when "11011" => level_vec_out <= "1111111111111111111011110111011111111111111111011110111011111111";
                    when "11100" => level_vec_out <= "1111111111111111111011110111011111111111111111111110111011111111";
                    when "11101" => level_vec_out <= "1111111111111111111011110111011111111111111111111110111011111111";
                    when "11110" => level_vec_out <= "1111111111111111111011110111111111111111111111111110111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111110111111111111111111111111110111111111111";
                when others => null;
                end case;
            when "011" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1011100100111111011000011011101101010110010000111101100000101101";
                    when "00001" => level_vec_out <= "1011100100111111011000011011101101010110010000111101100000101101";
                    when "00010" => level_vec_out <= "1011100100111111011000011011101101010110010000111101100000101101";
                    when "00011" => level_vec_out <= "1011100100111111011000011011101101010110010000111101100001101101";
                    when "00100" => level_vec_out <= "1011100100111111011100011011101101010110010000111101100001101101";
                    when "00101" => level_vec_out <= "1011100100111111011100011011101101010110010000111101100001101101";
                    when "00110" => level_vec_out <= "1011100101111111011100011011101101010110010000111101100001101101";
                    when "00111" => level_vec_out <= "1011100101111111011110011011101101010110010000111101100001101101";
                    when "01000" => level_vec_out <= "1011100101111111011110011011101101010110110000111101100001101111";
                    when "01001" => level_vec_out <= "1011100101111111011110011011101101110110110000111101100001101111";
                    when "01010" => level_vec_out <= "1011100101111111011110011011101101110110110000111101100001101111";
                    when "01011" => level_vec_out <= "1011110101111111011110011011101111110110110000111101100001101111";
                    when "01100" => level_vec_out <= "1011110101111111011110011011101111111110110000111101100001101111";
                    when "01101" => level_vec_out <= "1011110101111111011110011011101111111110110000111101100001111111";
                    when "01110" => level_vec_out <= "1011110101111111011110011011101111111110110000111101100001111111";
                    when "01111" => level_vec_out <= "1011110101111111011110011011101111111110110010111111100001111111";
                    when "10000" => level_vec_out <= "1011110101111111011110011011101111111110110010111111100001111111";
                    when "10001" => level_vec_out <= "1011110101111111111110011011101111111110111011111111100001111111";
                    when "10010" => level_vec_out <= "1011110101111111111110011011101111111110111011111111100011111111";
                    when "10011" => level_vec_out <= "1011110101111111111110011011101111111110111011111111100011111111";
                    when "10100" => level_vec_out <= "1111110111111111111110011011101111111110111011111111100011111111";
                    when "10101" => level_vec_out <= "1111110111111111111110011011101111111110111011111111100011111111";
                    when "10110" => level_vec_out <= "1111111111111111111110011011111111111110111011111111100011111111";
                    when "10111" => level_vec_out <= "1111111111111111111110011011111111111110111111111111100011111111";
                    when "11000" => level_vec_out <= "1111111111111111111110011011111111111110111111111111101011111111";
                    when "11001" => level_vec_out <= "1111111111111111111111011011111111111110111111111111101111111111";
                    when "11010" => level_vec_out <= "1111111111111111111111011111111111111110111111111111101111111111";
                    when "11011" => level_vec_out <= "1111111111111111111111011111111111111110111111111111101111111111";
                    when "11100" => level_vec_out <= "1111111111111111111111011111111111111110111111111111101111111111";
                    when "11101" => level_vec_out <= "1111111111111111111111111111111111111110111111111111101111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111110111111111111101111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111110111111111111101111111111";
                when others => null;
                end case;
            when "100" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1111110010101001001011010010110100101110110110110010010001000011";
                    when "00001" => level_vec_out <= "1111110010101001001011010010110100101110110110111010010001000011";
                    when "00010" => level_vec_out <= "1111110010101001001011010010110100101110110110111010010001000011";
                    when "00011" => level_vec_out <= "1111110010101001001011010010110100101110110110111010010001000011";
                    when "00100" => level_vec_out <= "1111110010101001001011010010110100101110110110111010010001000011";
                    when "00101" => level_vec_out <= "1111110010101011001011010010110100101110111110111010010001000011";
                    when "00110" => level_vec_out <= "1111110010101011001011010010110100101111111110111010010001000011";
                    when "00111" => level_vec_out <= "1111110010101011001011010010110100101111111110111010011001000011";
                    when "01000" => level_vec_out <= "1111110010111011001011010010110100101111111110111010011001000011";
                    when "01001" => level_vec_out <= "1111110010111011001011010010110100101111111110111010011001000011";
                    when "01010" => level_vec_out <= "1111110010111011001011010010111100101111111110111010011001000011";
                    when "01011" => level_vec_out <= "1111110010111011001011010010111100101111111110111010011001000111";
                    when "01100" => level_vec_out <= "1111110010111011001011010010111100101111111110111010011001000111";
                    when "01101" => level_vec_out <= "1111111010111111001011010010111100101111111110111010011001000111";
                    when "01110" => level_vec_out <= "1111111010111111001011010010111100111111111111111010011001000111";
                    when "01111" => level_vec_out <= "1111111010111111001011010010111100111111111111111010011001001111";
                    when "10000" => level_vec_out <= "1111111010111111001011010011111100111111111111111110011001001111";
                    when "10001" => level_vec_out <= "1111111010111111001011010011111100111111111111111110011011001111";
                    when "10010" => level_vec_out <= "1111111010111111001011010011111100111111111111111111011011001111";
                    when "10011" => level_vec_out <= "1111111010111111101111010011111110111111111111111111011011001111";
                    when "10100" => level_vec_out <= "1111111010111111101111010011111110111111111111111111011011001111";
                    when "10101" => level_vec_out <= "1111111010111111101111111011111110111111111111111111011011001111";
                    when "10110" => level_vec_out <= "1111111010111111101111111011111110111111111111111111011011001111";
                    when "10111" => level_vec_out <= "1111111010111111101111111011111110111111111111111111011111001111";
                    when "11000" => level_vec_out <= "1111111010111111101111111011111110111111111111111111011111101111";
                    when "11001" => level_vec_out <= "1111111010111111101111111011111110111111111111111111011111111111";
                    when "11010" => level_vec_out <= "1111111111111111111111111011111110111111111111111111011111111111";
                    when "11011" => level_vec_out <= "1111111111111111111111111011111110111111111111111111111111111111";
                    when "11100" => level_vec_out <= "1111111111111111111111111011111110111111111111111111111111111111";
                    when "11101" => level_vec_out <= "1111111111111111111111111011111111111111111111111111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111011111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "101" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0001101010100100101001011111101010010011011101111110011110000101";
                    when "00001" => level_vec_out <= "0001101010100100101001011111101010010111011101111110011110000101";
                    when "00010" => level_vec_out <= "0001101110100100101001011111101010010111011111111110011110000101";
                    when "00011" => level_vec_out <= "0001101110100100101001111111101010010111011111111110011110000101";
                    when "00100" => level_vec_out <= "0001101110100110101011111111101010010111011111111110011110000101";
                    when "00101" => level_vec_out <= "0001101110100110101011111111101010010111011111111110011110000101";
                    when "00110" => level_vec_out <= "0001101110100110101011111111101010010111011111111110011110100101";
                    when "00111" => level_vec_out <= "0001101110100110101011111111101010011111011111111110011110100101";
                    when "01000" => level_vec_out <= "0001101110101110101011111111101010011111011111111110011110100101";
                    when "01001" => level_vec_out <= "0001101110101111101011111111101010011111011111111110011110100101";
                    when "01010" => level_vec_out <= "0001101110101111101011111111101010011111011111111110011110101111";
                    when "01011" => level_vec_out <= "0001101110101111111011111111101010011111011111111110011110101111";
                    when "01100" => level_vec_out <= "0001101110101111111011111111101010011111011111111110011111101111";
                    when "01101" => level_vec_out <= "0011101110101111111011111111101010111111011111111110011111101111";
                    when "01110" => level_vec_out <= "0011101110101111111011111111101010111111011111111111011111101111";
                    when "01111" => level_vec_out <= "0111101110101111111011111111101010111111011111111111011111101111";
                    when "10000" => level_vec_out <= "0111101110101111111011111111101010111111011111111111011111101111";
                    when "10001" => level_vec_out <= "0111101110101111111011111111101010111111011111111111011111101111";
                    when "10010" => level_vec_out <= "0111101110111111111011111111101010111111111111111111011111101111";
                    when "10011" => level_vec_out <= "1111101110111111111011111111101010111111111111111111011111111111";
                    when "10100" => level_vec_out <= "1111101110111111111111111111101010111111111111111111011111111111";
                    when "10101" => level_vec_out <= "1111101110111111111111111111101010111111111111111111011111111111";
                    when "10110" => level_vec_out <= "1111101110111111111111111111101010111111111111111111111111111111";
                    when "10111" => level_vec_out <= "1111101111111111111111111111101010111111111111111111111111111111";
                    when "11000" => level_vec_out <= "1111101111111111111111111111101010111111111111111111111111111111";
                    when "11001" => level_vec_out <= "1111101111111111111111111111101010111111111111111111111111111111";
                    when "11010" => level_vec_out <= "1111101111111111111111111111101010111111111111111111111111111111";
                    when "11011" => level_vec_out <= "1111101111111111111111111111101011111111111111111111111111111111";
                    when "11100" => level_vec_out <= "1111101111111111111111111111111111111111111111111111111111111111";
                    when "11101" => level_vec_out <= "1111101111111111111111111111111111111111111111111111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "110" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0001100111010101011010110011001010011000001110110111110001101110";
                    when "00001" => level_vec_out <= "0001100111010101011010110111001010011000001110110111110001101110";
                    when "00010" => level_vec_out <= "0001110111010101011010110111001010011000001110110111110001101110";
                    when "00011" => level_vec_out <= "0001110111010101011010110111001010011010001110110111110001101110";
                    when "00100" => level_vec_out <= "0001110111010101011010110111001010011010001111110111111001101110";
                    when "00101" => level_vec_out <= "0001110111110101011010110111001010011010011111110111111001101110";
                    when "00110" => level_vec_out <= "1001110111110101011010110111001010011010011111110111111001101110";
                    when "00111" => level_vec_out <= "1001110111110101011010111111101010011010111111110111111001101110";
                    when "01000" => level_vec_out <= "1001110111110101011010111111101010011010111111110111111001101110";
                    when "01001" => level_vec_out <= "1001110111110101011010111111101010011010111111110111111101101110";
                    when "01010" => level_vec_out <= "1001110111110101111010111111101010011010111111110111111101101110";
                    when "01011" => level_vec_out <= "1001110111110101111010111111101110111010111111110111111101101110";
                    when "01100" => level_vec_out <= "1101110111110101111010111111101110111010111111110111111101101110";
                    when "01101" => level_vec_out <= "1101110111110101111010111111101110111010111111110111111101101110";
                    when "01110" => level_vec_out <= "1101110111110101111010111111101110111010111111110111111101111110";
                    when "01111" => level_vec_out <= "1101110111110101111010111111101111111010111111110111111101111110";
                    when "10000" => level_vec_out <= "1101110111110101111010111111101111111010111111110111111101111110";
                    when "10001" => level_vec_out <= "1101110111110101111010111111101111111010111111110111111101111110";
                    when "10010" => level_vec_out <= "1101110111110101111110111111101111111010111111110111111101111110";
                    when "10011" => level_vec_out <= "1101110111110101111110111111101111111010111111110111111101111110";
                    when "10100" => level_vec_out <= "1101110111110101111110111111101111111010111111110111111101111110";
                    when "10101" => level_vec_out <= "1101110111110101111111111111101111111011111111110111111101111110";
                    when "10110" => level_vec_out <= "1101110111110101111111111111101111111011111111110111111111111110";
                    when "10111" => level_vec_out <= "1101110111110101111111111111101111111011111111110111111111111110";
                    when "11000" => level_vec_out <= "1101110111110101111111111111101111111011111111111111111111111110";
                    when "11001" => level_vec_out <= "1101111111110101111111111111101111111011111111111111111111111110";
                    when "11010" => level_vec_out <= "1101111111110111111111111111101111111011111111111111111111111110";
                    when "11011" => level_vec_out <= "1101111111111111111111111111101111111011111111111111111111111110";
                    when "11100" => level_vec_out <= "1111111111111111111111111111101111111011111111111111111111111111";
                    when "11101" => level_vec_out <= "1111111111111111111111111111101111111011111111111111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111011111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111011111111111111111111111111";
                when others => null;
                end case;
            when "111" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1000100010011001100011110001010111001010000110000001000001110000";
                    when "00001" => level_vec_out <= "1000100010011001100011110011010111101010000110000101000001110000";
                    when "00010" => level_vec_out <= "1000100010011001100011110011010111101010000110000101000001110000";
                    when "00011" => level_vec_out <= "1000100010011001100011110011010111101010100110000101101001110000";
                    when "00100" => level_vec_out <= "1000100010011001100011110011010111101010100110000101101001110000";
                    when "00101" => level_vec_out <= "1000100011011001100011110011010111101010100110000101101001110000";
                    when "00110" => level_vec_out <= "1100100011011001100011110011010111101010100110000101101001110000";
                    when "00111" => level_vec_out <= "1100100011011001100011110011010111101010100110000101101001110000";
                    when "01000" => level_vec_out <= "1100100011011001100011110011010111101010100111000101101001110000";
                    when "01001" => level_vec_out <= "1100101011011001100011110011010111101010100111001101101001110000";
                    when "01010" => level_vec_out <= "1100101011011001100011110011010111101010101111001101101001110000";
                    when "01011" => level_vec_out <= "1100101011111001100011110011010111101010101111001101101001110000";
                    when "01100" => level_vec_out <= "1100111011111001100011110011010111101010101111001101101001110000";
                    when "01101" => level_vec_out <= "1100111011111001100011110011011111101010101111001111101001110000";
                    when "01110" => level_vec_out <= "1100111011111001100011111011011111101010101111001111101001110000";
                    when "01111" => level_vec_out <= "1100111011111001100011111011011111101010111111001111101001110000";
                    when "10000" => level_vec_out <= "1110111011111001100011111011011111101010111111001111101001111100";
                    when "10001" => level_vec_out <= "1110111011111001100011111011011111101010111111001111101001111100";
                    when "10010" => level_vec_out <= "1110111011111001100011111011011111101010111111001111101001111100";
                    when "10011" => level_vec_out <= "1111111011111001100011111011011111111010111111001111101001111100";
                    when "10100" => level_vec_out <= "1111111011111001100011111011011111111010111111001111101001111100";
                    when "10101" => level_vec_out <= "1111111011111001100011111011011111111010111111001111101001111100";
                    when "10110" => level_vec_out <= "1111111011111001100011111011011111111011111111011111101001111100";
                    when "10111" => level_vec_out <= "1111111011111001100011111011011111111111111111011111101001111100";
                    when "11000" => level_vec_out <= "1111111011111001100011111011011111111111111111111111111001111100";
                    when "11001" => level_vec_out <= "1111111011111001100011111011011111111111111111111111111001111100";
                    when "11010" => level_vec_out <= "1111111011111101100011111011011111111111111111111111111001111100";
                    when "11011" => level_vec_out <= "1111111011111101110011111011111111111111111111111111111001111100";
                    when "11100" => level_vec_out <= "1111111011111101111011111011111111111111111111111111111001111110";
                    when "11101" => level_vec_out <= "1111111011111101111011111011111111111111111111111111111011111110";
                    when "11110" => level_vec_out <= "1111111111111101111011111111111111111111111111111111111011111110";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111011111111";
                when others => null;
                end case;
            when others => null;
        end case;
    end process;
end Behavioral;