/**
 * @file level_hvec_gen_hdl.hpp
 * @brief This script generates HDL code for generating high-dimensional LEVEL vectors.
 * It is a novel method; for more information, please refer to our paper.
 *
 * @author Saeid Jamili and Marco Angioli
 * @note Author names are listed in alphabetical order.
 * @email <saeid.jamili@uniroma1.it>
 * @email <marco.angioli@uniroma1.it>
 *
 * @contributors
 *
 * @date Created: 24th July 2023
 * @date Last Updated: 23th August 2023
 *
 * @version 1.0.0
 *
 * @institute Sapienza University of Rome
 * @cite https://doi.org/10.xxxx/yyyyy
 *
 * @section DEPENDENCIES
 * - Dependency1: Description or version details.
 * - Dependency2: Description or version details.
 *
 * @section LICENSE
 * This file is part of the Aeneas HyperCompute Platform.
 *
 * Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 *
 * @section CHANGELOG
 * @version 1.0.0-dev - 23th August 2023
 * - Initial release
 *
 * @todo
 * - Complete level vector generator function
 * - Add training
 *
 * @see
 * -
 * -
 * -
 *
 */

module level_hvec_gen #(parameter int DI_PARALLEL_W_BITS = 64) (
  input logic [2:0] frame_index,
  input logic [4:0] frame_id,
  output logic [DI_PARALLEL_W_BITS-1:0] level_vec_out
);
  always_comb begin
    case (frame_index)
      0:
        case (frame_id)
          0:
            level_vec_out = 64'b0110110011110011111011100000011101101011001100000101111000100011;
          1:
            level_vec_out = 64'b0111110011110111111011100000011101101011001100000101111000100011;
          2:
            level_vec_out = 64'b0111110011110111111011100000011101101011001100000101111000100011;
          3:
            level_vec_out = 64'b0111110011110111111011100000011101101011001100100101111000100011;
          4:
            level_vec_out = 64'b0111110011110111111011100000011101101011001100100101111000100011;
          5:
            level_vec_out = 64'b0111110011110111111011100000011101101011001100100101111000100011;
          6:
            level_vec_out = 64'b0111110011110111111111100000011101101011001100100101111000100011;
          7:
            level_vec_out = 64'b0111110011110111111111100000011101101011011100100101111000100011;
          8:
            level_vec_out = 64'b0111110011111111111111100000011101101011011100100101111000100011;
          9:
            level_vec_out = 64'b0111110011111111111111100000011101101011011100100101111000100011;
          10:
            level_vec_out = 64'b0111110011111111111111100000011101101011111100100101111001100011;
          11:
            level_vec_out = 64'b0111111011111111111111100000011101101011111100101101111001100011;
          12:
            level_vec_out = 64'b0111111011111111111111100000011101101011111100101101111001100011;
          13:
            level_vec_out = 64'b0111111011111111111111100000011101101011111100101101111001100011;
          14:
            level_vec_out = 64'b0111111011111111111111100000011101101011111100111101111001100011;
          15:
            level_vec_out = 64'b0111111011111111111111100000011101101011111100111101111001100011;
          16:
            level_vec_out = 64'b0111111011111111111111101000011101101011111100111111111001100011;
          17:
            level_vec_out = 64'b0111111011111111111111101000011111101011111100111111111001100011;
          18:
            level_vec_out = 64'b0111111011111111111111101000011111101011111100111111111001101011;
          19:
            level_vec_out = 64'b0111111011111111111111101100011111101011111100111111111011101011;
          20:
            level_vec_out = 64'b0111111011111111111111101100011111101011111100111111111011111011;
          21:
            level_vec_out = 64'b0111111011111111111111101100011111101011111100111111111011111011;
          22:
            level_vec_out = 64'b0111111011111111111111101100011111101011111101111111111011111011;
          23:
            level_vec_out = 64'b0111111011111111111111101100011111101011111101111111111011111011;
          24:
            level_vec_out = 64'b0111111011111111111111101100011111111011111101111111111011111011;
          25:
            level_vec_out = 64'b0111111011111111111111111100011111111011111101111111111111111011;
          26:
            level_vec_out = 64'b0111111011111111111111111100011111111111111101111111111111111011;
          27:
            level_vec_out = 64'b1111111011111111111111111110011111111111111101111111111111111011;
          28:
            level_vec_out = 64'b1111111011111111111111111111011111111111111111111111111111111111;
          29:
            level_vec_out = 64'b1111111011111111111111111111011111111111111111111111111111111111;
          30:
            level_vec_out = 64'b1111111011111111111111111111011111111111111111111111111111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111011111111111111111111111111111111111;
        endcase
      1:
        case (frame_id)
          0:
            level_vec_out = 64'b1011001110101111000000000000010001001110000001001011000000101001;
          1:
            level_vec_out = 64'b1011001110101111000000000000010001001110000001001011100000101001;
          2:
            level_vec_out = 64'b1011001110101111000000000001010001101110000001001011100000101001;
          3:
            level_vec_out = 64'b1011001110101111100000000001010001111110000001011011100000101001;
          4:
            level_vec_out = 64'b1011001110101111100000000001010001111110000001111011100000101001;
          5:
            level_vec_out = 64'b1011001110101111100100100001010101111110000001111011100000101001;
          6:
            level_vec_out = 64'b1011001110101111100100100001010101111110000001111011100000101001;
          7:
            level_vec_out = 64'b1011001110101111100100100001110101111110000101111111100000101001;
          8:
            level_vec_out = 64'b1011001110101111100100100001110111111110000101111111100000101001;
          9:
            level_vec_out = 64'b1011001111101111100100100001110111111110001101111111100000101001;
          10:
            level_vec_out = 64'b1011011111101111100100100001110111111110001101111111100000101001;
          11:
            level_vec_out = 64'b1011011111101111100100100001110111111110001101111111100000101101;
          12:
            level_vec_out = 64'b1011011111101111100100100001110111111110001101111111100000101101;
          13:
            level_vec_out = 64'b1011011111101111100100100001110111111110001101111111101001101101;
          14:
            level_vec_out = 64'b1011011111101111100100100001110111111110001101111111101001101101;
          15:
            level_vec_out = 64'b1011011111111111100100100001110111111110001101111111101001101101;
          16:
            level_vec_out = 64'b1011011111111111100100100011110111111110001101111111101011101101;
          17:
            level_vec_out = 64'b1011011111111111100100101011110111111110101111111111101011101101;
          18:
            level_vec_out = 64'b1011011111111111100100101011110111111110111111111111101011101101;
          19:
            level_vec_out = 64'b1011011111111111110100101011110111111110111111111111101011101101;
          20:
            level_vec_out = 64'b1011011111111111110100101011110111111110111111111111101111101101;
          21:
            level_vec_out = 64'b1011111111111111110100111111110111111110111111111111101111101101;
          22:
            level_vec_out = 64'b1011111111111111110101111111110111111110111111111111101111101111;
          23:
            level_vec_out = 64'b1111111111111111110101111111110111111110111111111111101111101111;
          24:
            level_vec_out = 64'b1111111111111111110101111111110111111110111111111111101111101111;
          25:
            level_vec_out = 64'b1111111111111111110101111111110111111111111111111111101111101111;
          26:
            level_vec_out = 64'b1111111111111111110101111111110111111111111111111111101111101111;
          27:
            level_vec_out = 64'b1111111111111111110111111111110111111111111111111111101111101111;
          28:
            level_vec_out = 64'b1111111111111111110111111111110111111111111111111111101111101111;
          29:
            level_vec_out = 64'b1111111111111111110111111111110111111111111111111111101111101111;
          30:
            level_vec_out = 64'b1111111111111111111111111111110111111111111111111111101111101111;
          31:
            level_vec_out = 64'b1111111111111111111111111111110111111111111111111111111111101111;
        endcase
      2:
        case (frame_id)
          0:
            level_vec_out = 64'b1111100000101111101110001110110100110100010110011111101011011010;
          1:
            level_vec_out = 64'b1111101000101111101110001110110100110100010110011111101011011010;
          2:
            level_vec_out = 64'b1111101000101111101110001110110100110100010110011111101011011010;
          3:
            level_vec_out = 64'b1111101000101111101110001110110100110100010110011111101011111010;
          4:
            level_vec_out = 64'b1111101000101111101110001110110100110100010110011111101011111010;
          5:
            level_vec_out = 64'b1111101000101111101110001110110110110100010111011111101011111010;
          6:
            level_vec_out = 64'b1111101001101111101110001110110110110100010111011111101011111110;
          7:
            level_vec_out = 64'b1111101001101111101110001110110110111100010111011111101011111110;
          8:
            level_vec_out = 64'b1111101001101111101110011110110110111100010111011111101011111110;
          9:
            level_vec_out = 64'b1111101001101111101110111110110110111100010111011111101011111110;
          10:
            level_vec_out = 64'b1111101001111111101111111110110110111100010111011111101011111110;
          11:
            level_vec_out = 64'b1111101001111111101111111110110110111100010111011111101011111110;
          12:
            level_vec_out = 64'b1111101101111111101111111110110110111100010111011111101111111110;
          13:
            level_vec_out = 64'b1111101101111111101111111110110110111100010111011111101111111110;
          14:
            level_vec_out = 64'b1111101101111111101111111110110110111100010111011111101111111110;
          15:
            level_vec_out = 64'b1111101101111111101111111110110110111100010111111111101111111110;
          16:
            level_vec_out = 64'b1111101101111111101111111110110110111100010111111111101111111110;
          17:
            level_vec_out = 64'b1111101101111111101111111110110110111100010111111111101111111110;
          18:
            level_vec_out = 64'b1111101101111111101111111110110110111100110111111111101111111110;
          19:
            level_vec_out = 64'b1111101101111111101111111110110110111100111111111111101111111110;
          20:
            level_vec_out = 64'b1111101111111111101111111110110110111100111111111111101111111110;
          21:
            level_vec_out = 64'b1111111111111111101111111110110110111101111111111111101111111110;
          22:
            level_vec_out = 64'b1111111111111111101111111110110110111111111111111111101111111110;
          23:
            level_vec_out = 64'b1111111111111111101111111111110110111111111111111111101111111110;
          24:
            level_vec_out = 64'b1111111111111111101111111111110110111111111111111111101111111110;
          25:
            level_vec_out = 64'b1111111111111111101111111111110110111111111111111111101111111110;
          26:
            level_vec_out = 64'b1111111111111111111111111111110111111111111111111111101111111110;
          27:
            level_vec_out = 64'b1111111111111111111111111111110111111111111111111111101111111110;
          28:
            level_vec_out = 64'b1111111111111111111111111111110111111111111111111111111111111110;
          29:
            level_vec_out = 64'b1111111111111111111111111111110111111111111111111111111111111110;
          30:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111110;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        endcase
      3:
        case (frame_id)
          0:
            level_vec_out = 64'b1111100100011001001101101111101001101101111000011011110111111001;
          1:
            level_vec_out = 64'b1111101100011001001101101111101001101101111000011011110111111001;
          2:
            level_vec_out = 64'b1111101100011001001101101111101001101101111000011011110111111001;
          3:
            level_vec_out = 64'b1111101100011001001101101111101001101101111000011011110111111001;
          4:
            level_vec_out = 64'b1111101100011001001101101111101011101101111000011011110111111001;
          5:
            level_vec_out = 64'b1111101100011001001101101111101011101101111000011011110111111001;
          6:
            level_vec_out = 64'b1111101100011001001101101111101011101101111000011011110111111001;
          7:
            level_vec_out = 64'b1111101100011001001101101111101011101101111000011011110111111001;
          8:
            level_vec_out = 64'b1111101101011001001101101111101011101101111000011011110111111001;
          9:
            level_vec_out = 64'b1111101101011001001101101111101011101111111000111011111111111001;
          10:
            level_vec_out = 64'b1111101101011001001101101111101011101111111000111011111111111001;
          11:
            level_vec_out = 64'b1111101101011001001101101111101011101111111000111011111111111001;
          12:
            level_vec_out = 64'b1111101101011001001101101111101011101111111000111011111111111001;
          13:
            level_vec_out = 64'b1111101101011001001101101111101011101111111001111011111111111001;
          14:
            level_vec_out = 64'b1111101101011001001101101111101011111111111001111011111111111001;
          15:
            level_vec_out = 64'b1111101101011001001101101111101011111111111001111011111111111001;
          16:
            level_vec_out = 64'b1111101101011001001101101111101011111111111001111011111111111001;
          17:
            level_vec_out = 64'b1111101101011001001101101111101111111111111001111011111111111001;
          18:
            level_vec_out = 64'b1111101101011001001101111111101111111111111001111011111111111001;
          19:
            level_vec_out = 64'b1111101101011101001101111111101111111111111001111011111111111001;
          20:
            level_vec_out = 64'b1111101101111101001101111111101111111111111001111011111111111001;
          21:
            level_vec_out = 64'b1111101101111101001101111111101111111111111001111011111111111001;
          22:
            level_vec_out = 64'b1111101101111101001101111111101111111111111001111011111111111001;
          23:
            level_vec_out = 64'b1111101101111101001111111111101111111111111001111011111111111001;
          24:
            level_vec_out = 64'b1111101101111101001111111111111111111111111001111011111111111101;
          25:
            level_vec_out = 64'b1111101101111101001111111111111111111111111101111011111111111101;
          26:
            level_vec_out = 64'b1111101101111101011111111111111111111111111101111011111111111101;
          27:
            level_vec_out = 64'b1111101101111101011111111111111111111111111101111011111111111101;
          28:
            level_vec_out = 64'b1111101101111101011111111111111111111111111101111011111111111111;
          29:
            level_vec_out = 64'b1111111101111101011111111111111111111111111101111111111111111111;
          30:
            level_vec_out = 64'b1111111111111101011111111111111111111111111111111111111111111111;
          31:
            level_vec_out = 64'b1111111111111101011111111111111111111111111111111111111111111111;
        endcase
      4:
        case (frame_id)
          0:
            level_vec_out = 64'b0111110011111110101011011101010011001001011110110111000001000011;
          1:
            level_vec_out = 64'b0111110011111110101011011101010011001001011111110111000001000011;
          2:
            level_vec_out = 64'b0111110011111110101011011101010011001001011111110111000001001011;
          3:
            level_vec_out = 64'b0111110011111110101011011101010011001001011111110111000001001011;
          4:
            level_vec_out = 64'b0111110011111110101011011111010011011001011111110111010001001011;
          5:
            level_vec_out = 64'b0111110011111111101011011111010011011001011111110111010001001011;
          6:
            level_vec_out = 64'b0111110011111111101011011111010011011001011111110111010001001011;
          7:
            level_vec_out = 64'b0111110011111111101011011111010011011001011111110111010001001011;
          8:
            level_vec_out = 64'b0111110011111111101011011111010011011001011111110111010001001011;
          9:
            level_vec_out = 64'b0111110011111111101011011111010011011001011111110111010001001011;
          10:
            level_vec_out = 64'b0111110011111111101011011111010011011001011111110111010001001011;
          11:
            level_vec_out = 64'b0111110011111111111011011111010011011001011111111111010001001011;
          12:
            level_vec_out = 64'b0111110011111111111011011111010011011001011111111111011001001011;
          13:
            level_vec_out = 64'b0111110011111111111011011111010011011001011111111111011001001011;
          14:
            level_vec_out = 64'b0111110011111111111011011111010011011001011111111111011001001011;
          15:
            level_vec_out = 64'b0111110011111111111011111111010011011001011111111111011001001011;
          16:
            level_vec_out = 64'b0111110011111111111011111111010011111101011111111111011001001011;
          17:
            level_vec_out = 64'b0111110111111111111011111111010011111101011111111111011001001011;
          18:
            level_vec_out = 64'b0111110111111111111011111111010011111101011111111111011001001111;
          19:
            level_vec_out = 64'b0111110111111111111011111111010011111101011111111111011001001111;
          20:
            level_vec_out = 64'b0111110111111111111011111111010011111101011111111111011001001111;
          21:
            level_vec_out = 64'b0111110111111111111011111111011011111111011111111111011001001111;
          22:
            level_vec_out = 64'b0111110111111111111011111111011011111111011111111111011001001111;
          23:
            level_vec_out = 64'b0111110111111111111011111111011011111111011111111111011011101111;
          24:
            level_vec_out = 64'b1111111111111111111011111111111011111111011111111111011011101111;
          25:
            level_vec_out = 64'b1111111111111111111011111111111011111111011111111111011011101111;
          26:
            level_vec_out = 64'b1111111111111111111011111111111011111111011111111111011011111111;
          27:
            level_vec_out = 64'b1111111111111111111011111111111011111111011111111111111111111111;
          28:
            level_vec_out = 64'b1111111111111111111011111111111011111111011111111111111111111111;
          29:
            level_vec_out = 64'b1111111111111111111111111111111011111111111111111111111111111111;
          30:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        endcase
      5:
        case (frame_id)
          0:
            level_vec_out = 64'b1001000100000001110110111101010001111000001001100010001000010110;
          1:
            level_vec_out = 64'b1001000100000001110110111101010001111000001001100010001000010110;
          2:
            level_vec_out = 64'b1001000100000001110110111101010011111000001001100010001100011110;
          3:
            level_vec_out = 64'b1001000100000001110110111101010011111000001001100010001100011110;
          4:
            level_vec_out = 64'b1001000100000001110110111101010011111000001001100010001100011110;
          5:
            level_vec_out = 64'b1001000100000001110110111101010011111000001001100010001100011111;
          6:
            level_vec_out = 64'b1001000100000001110110111101010011111000001001101010001100011111;
          7:
            level_vec_out = 64'b1001000110100001110110111101010011111000001001101010001100011111;
          8:
            level_vec_out = 64'b1001001110100001110110111101010011111000001001101010001100011111;
          9:
            level_vec_out = 64'b1001001110100001110110111101010011111000001001101010001100011111;
          10:
            level_vec_out = 64'b1001001110100001110110111101010011111000001001101010001100011111;
          11:
            level_vec_out = 64'b1001001110100001110110111111010011111000001001101010001100011111;
          12:
            level_vec_out = 64'b1101011110100001110110111111010011111000011001111010101100011111;
          13:
            level_vec_out = 64'b1111011110100001110110111111010111111000011001111010101110011111;
          14:
            level_vec_out = 64'b1111011110100001110110111111010111111000011001111110101110011111;
          15:
            level_vec_out = 64'b1111011110100001110111111111010111111000011001111111101110011111;
          16:
            level_vec_out = 64'b1111011110100001110111111111010111111000011001111111101110011111;
          17:
            level_vec_out = 64'b1111011110100001110111111111010111111000011001111111101110011111;
          18:
            level_vec_out = 64'b1111011110100001110111111111010111111000011101111111111110011111;
          19:
            level_vec_out = 64'b1111011111100101110111111111010111111000011101111111111110011111;
          20:
            level_vec_out = 64'b1111011111101101110111111111010111111010011101111111111110011111;
          21:
            level_vec_out = 64'b1111011111101101110111111111011111111010011101111111111110011111;
          22:
            level_vec_out = 64'b1111011111101101110111111111011111111010011101111111111110011111;
          23:
            level_vec_out = 64'b1111011111101101110111111111011111111010011101111111111110111111;
          24:
            level_vec_out = 64'b1111011111101101110111111111011111111010011101111111111110111111;
          25:
            level_vec_out = 64'b1111011111101111110111111111011111111010011101111111111110111111;
          26:
            level_vec_out = 64'b1111011111101111110111111111011111111010011101111111111111111111;
          27:
            level_vec_out = 64'b1111011111101111110111111111011111111010011111111111111111111111;
          28:
            level_vec_out = 64'b1111111111101111110111111111011111111010011111111111111111111111;
          29:
            level_vec_out = 64'b1111111111101111110111111111011111111011011111111111111111111111;
          30:
            level_vec_out = 64'b1111111111101111110111111111011111111011011111111111111111111111;
          31:
            level_vec_out = 64'b1111111111111111110111111111111111111111111111111111111111111111;
        endcase
      6:
        case (frame_id)
          0:
            level_vec_out = 64'b0001101000011100100111001010110101101101011110000101010001001000;
          1:
            level_vec_out = 64'b0001101000011100100111001010110101101101011110000111010001001000;
          2:
            level_vec_out = 64'b0001101000011100100111001010110101101101011110000111010001001000;
          3:
            level_vec_out = 64'b0001101000011100110111001011110101101101011110000111010001001000;
          4:
            level_vec_out = 64'b0001101000011100110111001011110101101101011110000111010001001000;
          5:
            level_vec_out = 64'b0001101000011100110111001011110101101101011110000111010001001000;
          6:
            level_vec_out = 64'b0001101001011100110111001011111101111101011110000111010001001000;
          7:
            level_vec_out = 64'b0001101001011100110111001011111101111101011110100111010001001000;
          8:
            level_vec_out = 64'b0001101001011100110111001011111111111101011110100111010001001000;
          9:
            level_vec_out = 64'b0001101001011100110111001011111111111101011110100111010001001000;
          10:
            level_vec_out = 64'b0001101001011100110111001011111111111101011110100111010001001000;
          11:
            level_vec_out = 64'b0001101001011100110111001011111111111101011110100111010001001001;
          12:
            level_vec_out = 64'b0001101001011100110111001011111111111101011110100111010001001001;
          13:
            level_vec_out = 64'b0001101001011101110111001011111111111101011110100111010001001001;
          14:
            level_vec_out = 64'b0111101001011101110111001011111111111101011110101111010101001001;
          15:
            level_vec_out = 64'b0111101001011101110111001011111111111101011110101111010101011001;
          16:
            level_vec_out = 64'b0111101001011101110111001011111111111101011110111111010101011001;
          17:
            level_vec_out = 64'b0111101001011101110111011011111111111101011110111111010101011001;
          18:
            level_vec_out = 64'b0111101001011101110111011011111111111101011110111111010101011001;
          19:
            level_vec_out = 64'b0111101001011101110111011011111111111101011110111111010101011001;
          20:
            level_vec_out = 64'b1111101101011101110111011011111111111101011110111111010101011001;
          21:
            level_vec_out = 64'b1111101101011101110111011011111111111101011110111111010101011001;
          22:
            level_vec_out = 64'b1111101101011101111111011011111111111101011110111111010111011001;
          23:
            level_vec_out = 64'b1111111101011101111111011011111111111101011110111111011111011001;
          24:
            level_vec_out = 64'b1111111101011101111111011011111111111101011110111111011111011001;
          25:
            level_vec_out = 64'b1111111101011111111111011011111111111101011110111111011111011101;
          26:
            level_vec_out = 64'b1111111111011111111111011011111111111101011110111111011111011101;
          27:
            level_vec_out = 64'b1111111111011111111111011111111111111101011110111111011111011101;
          28:
            level_vec_out = 64'b1111111111011111111111011111111111111101111110111111111111011101;
          29:
            level_vec_out = 64'b1111111111011111111111011111111111111101111110111111111111111101;
          30:
            level_vec_out = 64'b1111111111011111111111111111111111111101111110111111111111111111;
          31:
            level_vec_out = 64'b1111111111011111111111111111111111111111111110111111111111111111;
        endcase
      7:
        case (frame_id)
          0:
            level_vec_out = 64'b1100010000101000011100110100100110101100101111101100000100010110;
          1:
            level_vec_out = 64'b1101010000101000011100110100100110101100101111101100000100010110;
          2:
            level_vec_out = 64'b1101010000101000011100110100100110101100101111101100100100010111;
          3:
            level_vec_out = 64'b1101010000101000011100110101100110101100101111101100100100010111;
          4:
            level_vec_out = 64'b1101011000101000111100110101101110101100101111101100100100010111;
          5:
            level_vec_out = 64'b1101011000101100111100110101101110101100101111101100100100010111;
          6:
            level_vec_out = 64'b1101011000101100111100110101101110101100101111101110100100010111;
          7:
            level_vec_out = 64'b1101011000101100111100110101101110101100101111101110100100010111;
          8:
            level_vec_out = 64'b1101011000101100111100110101101111101100101111101110101100010111;
          9:
            level_vec_out = 64'b1101011001101100111100110101101111101100101111111110101100010111;
          10:
            level_vec_out = 64'b1101011111101100111100110101101111101100101111111111101100010111;
          11:
            level_vec_out = 64'b1101011111101100111100110101101111101100101111111111101110010111;
          12:
            level_vec_out = 64'b1101011111101100111100110101101111101100101111111111101110010111;
          13:
            level_vec_out = 64'b1101011111101101111100110101101111101100101111111111101110010111;
          14:
            level_vec_out = 64'b1111011111101101111100110101101111101100101111111111101110010111;
          15:
            level_vec_out = 64'b1111011111101111111100110101101111101100101111111111101110110111;
          16:
            level_vec_out = 64'b1111011111101111111100110101101111111100101111111111101110110111;
          17:
            level_vec_out = 64'b1111011111101111111100110101101111111100101111111111101111110111;
          18:
            level_vec_out = 64'b1111011111101111111100110101101111111100111111111111101111110111;
          19:
            level_vec_out = 64'b1111011111101111111110110101101111111100111111111111101111110111;
          20:
            level_vec_out = 64'b1111011111101111111110110101101111111100111111111111101111110111;
          21:
            level_vec_out = 64'b1111011111101111111110110101101111111100111111111111101111110111;
          22:
            level_vec_out = 64'b1111111111101111111110110101101111111101111111111111101111110111;
          23:
            level_vec_out = 64'b1111111111101111111110110101101111111101111111111111101111110111;
          24:
            level_vec_out = 64'b1111111111101111111110110101111111111101111111111111111111110111;
          25:
            level_vec_out = 64'b1111111111101111111110110101111111111101111111111111111111111111;
          26:
            level_vec_out = 64'b1111111111101111111111110101111111111101111111111111111111111111;
          27:
            level_vec_out = 64'b1111111111111111111111110101111111111101111111111111111111111111;
          28:
            level_vec_out = 64'b1111111111111111111111110101111111111101111111111111111111111111;
          29:
            level_vec_out = 64'b1111111111111111111111110111111111111111111111111111111111111111;
          30:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        endcase
    endcase
  end
endmodule