----
 -- @file level_hvec_gen_hdl.hpp
 -- @brief This script generates HDL code for generating high-dimensional LEVEL vectors.
 -- It is a novel method; for more information, please refer to our paper.
 --
 -- @author Saeid Jamili and Marco Angioli
 -- @note Author names are listed in alphabetical order.
 -- @email <saeid.jamili@uniroma1.it>
 -- @email <marco.angioli@uniroma1.it>
 --
 -- @contributors
 --
 -- @date Created: 24th July 2023
 -- @date Last Updated: 23th August 2023
 --
 -- @version 1.0.0
 --
 -- @institute Sapienza University of Rome
 -- @cite https://doi.org/10.xxxx/yyyyy
 --
 -- @section DEPENDENCIES
 -- - Dependency1: Description or version details.
 -- - Dependency2: Description or version details.
 --
 -- @section LICENSE
 -- This file is part of the Aeneas HyperCompute Platform.
 --
 -- Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 --
 -- @section CHANGELOG
 -- @version 1.0.0-dev - 23th August 2023
 -- - Initial release
 --
 -- @todo
 -- - Complete level vector generator function
 -- - Add training
 --
 -- @see
 -- -
 -- -
 -- -
 --
 --

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity level_vec_gen is
    Port ( level_vec_out : out  STD_LOGIC_VECTOR (63 downto 0);
           frame_index : in  STD_LOGIC_VECTOR (2 downto 0);
           frame_id : in  STD_LOGIC_VECTOR (4 downto 0));
end level_vec_gen;

architecture Behavioral of level_vec_gen is
begin
    process (frame_index, frame_id)
    begin
        -- Update this function to match your requirements
        case frame_index is
            when "000" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1100111111011010111110111111110001101110110100000001100111100101";
                    when "00001" => level_vec_out <= "1100111111011010111110111111110001101110110100000001100111100101";
                    when "00010" => level_vec_out <= "1100111111011010111110111111111001101110110110000001100111100101";
                    when "00011" => level_vec_out <= "1100111111011010111110111111111001101110110110010001100111100101";
                    when "00100" => level_vec_out <= "1100111111011010111110111111111101101110110110010001100111100101";
                    when "00101" => level_vec_out <= "1100111111011010111110111111111101101110110110011001100111100101";
                    when "00110" => level_vec_out <= "1100111111011010111110111111111101101110110110011001101111100101";
                    when "00111" => level_vec_out <= "1100111111011010111110111111111101101110110110011001101111100101";
                    when "01000" => level_vec_out <= "1100111111011010111110111111111101101110110110011001101111100101";
                    when "01001" => level_vec_out <= "1111111111011010111110111111111101101110110110011001101111100101";
                    when "01010" => level_vec_out <= "1111111111011010111110111111111101101110110110011001101111100101";
                    when "01011" => level_vec_out <= "1111111111011010111110111111111101101110110110011001101111100101";
                    when "01100" => level_vec_out <= "1111111111011010111110111111111101111110110110011001101111100101";
                    when "01101" => level_vec_out <= "1111111111011010111110111111111111111110110110011001101111100101";
                    when "01110" => level_vec_out <= "1111111111011010111110111111111111111110110110011001101111100101";
                    when "01111" => level_vec_out <= "1111111111011010111110111111111111111110110110011001101111100101";
                    when "10000" => level_vec_out <= "1111111111011010111110111111111111111110110110011011101111100101";
                    when "10001" => level_vec_out <= "1111111111011010111110111111111111111110111110011011101111100101";
                    when "10010" => level_vec_out <= "1111111111011010111110111111111111111110111110011011101111100111";
                    when "10011" => level_vec_out <= "1111111111011010111110111111111111111110111110011011101111100111";
                    when "10100" => level_vec_out <= "1111111111011010111110111111111111111110111110011011101111100111";
                    when "10101" => level_vec_out <= "1111111111011010111110111111111111111110111110011011101111100111";
                    when "10110" => level_vec_out <= "1111111111111010111110111111111111111110111111111111101111100111";
                    when "10111" => level_vec_out <= "1111111111111010111110111111111111111110111111111111101111100111";
                    when "11000" => level_vec_out <= "1111111111111010111110111111111111111110111111111111101111100111";
                    when "11001" => level_vec_out <= "1111111111111010111110111111111111111110111111111111101111101111";
                    when "11010" => level_vec_out <= "1111111111111110111111111111111111111111111111111111101111101111";
                    when "11011" => level_vec_out <= "1111111111111110111111111111111111111111111111111111101111101111";
                    when "11100" => level_vec_out <= "1111111111111110111111111111111111111111111111111111101111101111";
                    when "11101" => level_vec_out <= "1111111111111110111111111111111111111111111111111111101111101111";
                    when "11110" => level_vec_out <= "1111111111111110111111111111111111111111111111111111111111101111";
                    when "11111" => level_vec_out <= "1111111111111110111111111111111111111111111111111111111111101111";
                when others => null;
                end case;
            when "001" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1100011000111011100010011001100010000000100110010110000011010010";
                    when "00001" => level_vec_out <= "1100011000111011100010011001100010000000100110010110000011010010";
                    when "00010" => level_vec_out <= "1100011000111011100010011001100010000010100110010110000011010010";
                    when "00011" => level_vec_out <= "1100011000111011100010011001100010000010100110010110000011010010";
                    when "00100" => level_vec_out <= "1100011000111011100010011101100010000010100110010110100011010010";
                    when "00101" => level_vec_out <= "1100011000111011100010011101100010000010100110010111100011010010";
                    when "00110" => level_vec_out <= "1100011000111011100010011101100010000010100110010111100011010010";
                    when "00111" => level_vec_out <= "1100011000111011100010011101100010000011100110010111100011010010";
                    when "01000" => level_vec_out <= "1100011000111011100010011101100010000011100110010111100011110010";
                    when "01001" => level_vec_out <= "1100011000111011100010011101110010000011100110010111100011110010";
                    when "01010" => level_vec_out <= "1100011000111011100010011101110010000011100110010111100011110010";
                    when "01011" => level_vec_out <= "1100011000111011100010011101110010000011110110110111100011110110";
                    when "01100" => level_vec_out <= "1100011000111011100010011101110010000011110110110111100011110110";
                    when "01101" => level_vec_out <= "1110011000111011100010011101110010000011110110110111100011110110";
                    when "01110" => level_vec_out <= "1110011000111011100010011101110010000011110110110111100011110110";
                    when "01111" => level_vec_out <= "1110011000111011100010011101110010100011110110110111100011110111";
                    when "10000" => level_vec_out <= "1110011000111011100010011101110010100011110110110111100011110111";
                    when "10001" => level_vec_out <= "1110011100111011100010011101110010100011110110110111100011110111";
                    when "10010" => level_vec_out <= "1110011100111011100010011101110010100011110111110111100011110111";
                    when "10011" => level_vec_out <= "1110011100111011100010011101110011100011110111110111101011110111";
                    when "10100" => level_vec_out <= "1110011100111011100010011111110011100011110111111111101011110111";
                    when "10101" => level_vec_out <= "1110011101111011100010011111110011100011110111111111111011110111";
                    when "10110" => level_vec_out <= "1110011101111011100010011111110011100011110111111111111011110111";
                    when "10111" => level_vec_out <= "1110011101111011100010011111110011100011110111111111111011110111";
                    when "11000" => level_vec_out <= "1110011101111011100010011111110011100111111111111111111011110111";
                    when "11001" => level_vec_out <= "1110011101111011100010011111110111100111111111111111111011110111";
                    when "11010" => level_vec_out <= "1110011101111011100010011111110111101111111111111111111011110111";
                    when "11011" => level_vec_out <= "1110011101111011100011011111110111101111111111111111111011110111";
                    when "11100" => level_vec_out <= "1110011101111111101111111111110111101111111111111111111011111111";
                    when "11101" => level_vec_out <= "1111011101111111101111111111110111101111111111111111111011111111";
                    when "11110" => level_vec_out <= "1111111101111111111111111111111111101111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "010" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1101000011100001101001010111100001100100010001011011010011101110";
                    when "00001" => level_vec_out <= "1101000011100001101001010111100001100100010001011011010011101110";
                    when "00010" => level_vec_out <= "1101000011100001101001010111100001100100010001011011010011111110";
                    when "00011" => level_vec_out <= "1101000011100001111001010111100001100100010001011011010011111110";
                    when "00100" => level_vec_out <= "1101000011100001111001010111100001100100010011011011010011111110";
                    when "00101" => level_vec_out <= "1101000011100001111001010111100001100100010011011011010011111110";
                    when "00110" => level_vec_out <= "1101000011100001111001010111100001100100010011011011010011111110";
                    when "00111" => level_vec_out <= "1101000011100001111001010111100001100100010011011011010011111110";
                    when "01000" => level_vec_out <= "1101000011100001111001010111100001100110010011011011010011111110";
                    when "01001" => level_vec_out <= "1101010011100001111001010111100001100110010011011011010011111110";
                    when "01010" => level_vec_out <= "1101010011100001111001010111100001110111010011011011010011111110";
                    when "01011" => level_vec_out <= "1101010011100001111001110111100001110111010011011011010011111110";
                    when "01100" => level_vec_out <= "1101011011100101111001110111100001110111010011111011010011111110";
                    when "01101" => level_vec_out <= "1101011011100101111001110111100011110111010011111011010011111110";
                    when "01110" => level_vec_out <= "1101011011100101111001110111100011110111010011111011010011111111";
                    when "01111" => level_vec_out <= "1101011011100101111001110111100011110111010011111111010011111111";
                    when "10000" => level_vec_out <= "1101011011100101111001110111100011111111010011111111010011111111";
                    when "10001" => level_vec_out <= "1101011111100101111001110111101011111111010011111111010011111111";
                    when "10010" => level_vec_out <= "1101011111100101111101110111101011111111010011111111010011111111";
                    when "10011" => level_vec_out <= "1101011111100101111111111111101011111111010011111111010011111111";
                    when "10100" => level_vec_out <= "1101011111100101111111111111101011111111010011111111010011111111";
                    when "10101" => level_vec_out <= "1101011111100101111111111111101011111111011011111111010011111111";
                    when "10110" => level_vec_out <= "1101011111100101111111111111101011111111011011111111010011111111";
                    when "10111" => level_vec_out <= "1101011111100101111111111111111011111111011011111111010011111111";
                    when "11000" => level_vec_out <= "1101111111100101111111111111111011111111011011111111011011111111";
                    when "11001" => level_vec_out <= "1101111111100101111111111111111111111111011011111111011011111111";
                    when "11010" => level_vec_out <= "1101111111100101111111111111111111111111011011111111111011111111";
                    when "11011" => level_vec_out <= "1101111111110101111111111111111111111111111011111111111011111111";
                    when "11100" => level_vec_out <= "1101111111110101111111111111111111111111111011111111111011111111";
                    when "11101" => level_vec_out <= "1101111111110101111111111111111111111111111111111111111011111111";
                    when "11110" => level_vec_out <= "1101111111110101111111111111111111111111111111111111111011111111";
                    when "11111" => level_vec_out <= "1111111111111101111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "011" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0111110001001110101001000111100111000101101010000101100111110101";
                    when "00001" => level_vec_out <= "0111110101001110101001000111101111000101101010000101100111111101";
                    when "00010" => level_vec_out <= "0111110101001110101001000111101111000101101010000101100111111101";
                    when "00011" => level_vec_out <= "0111110101001110101001000111101111000101101010000101100111111101";
                    when "00100" => level_vec_out <= "0111110101001110101001000111101111000111111010000101100111111101";
                    when "00101" => level_vec_out <= "0111110101001110101001000111101111000111111010000101100111111101";
                    when "00110" => level_vec_out <= "0111110101001110101001000111101111000111111010000101100111111111";
                    when "00111" => level_vec_out <= "0111110101001110101011000111101111000111111010000111100111111111";
                    when "01000" => level_vec_out <= "0111110101001110101011000111101111000111111010000111100111111111";
                    when "01001" => level_vec_out <= "0111110101001110101011010111101111000111111010000111100111111111";
                    when "01010" => level_vec_out <= "0111110101001110101011010111101111000111111010000111101111111111";
                    when "01011" => level_vec_out <= "0111110101001110101011010111101111000111111010000111101111111111";
                    when "01100" => level_vec_out <= "0111110101001110101011010111101111000111111010000111101111111111";
                    when "01101" => level_vec_out <= "0111110101001110101011010111111111000111111010000111101111111111";
                    when "01110" => level_vec_out <= "0111110101001110101011010111111111100111111110000111101111111111";
                    when "01111" => level_vec_out <= "0111110101001110101011010111111111100111111110100111101111111111";
                    when "10000" => level_vec_out <= "0111110101001110101011010111111111100111111110100111101111111111";
                    when "10001" => level_vec_out <= "0111110111001110101011011111111111100111111110100111101111111111";
                    when "10010" => level_vec_out <= "0111110111001110111011011111111111100111111110110111101111111111";
                    when "10011" => level_vec_out <= "0111110111001110111011011111111111100111111110110111101111111111";
                    when "10100" => level_vec_out <= "0111110111011110111011011111111111100111111110110111101111111111";
                    when "10101" => level_vec_out <= "0111110111011110111011011111111111100111111110110111101111111111";
                    when "10110" => level_vec_out <= "1111110111011110111011011111111111100111111110110111101111111111";
                    when "10111" => level_vec_out <= "1111110111011110111111011111111111100111111110110111101111111111";
                    when "11000" => level_vec_out <= "1111110111011110111111011111111111110111111110110111101111111111";
                    when "11001" => level_vec_out <= "1111110111011111111111011111111111110111111110110111101111111111";
                    when "11010" => level_vec_out <= "1111110111011111111111011111111111110111111110110111101111111111";
                    when "11011" => level_vec_out <= "1111110111011111111111111111111111110111111110111111101111111111";
                    when "11100" => level_vec_out <= "1111110111011111111111111111111111110111111110111111101111111111";
                    when "11101" => level_vec_out <= "1111110111011111111111111111111111111111111110111111111111111111";
                    when "11110" => level_vec_out <= "1111110111011111111111111111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111011111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "100" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1011101111001001001011101110001101100100001100110001110010101011";
                    when "00001" => level_vec_out <= "1011101111001001001011101110001101100100001100110001110010101011";
                    when "00010" => level_vec_out <= "1011101111001001101011101110001101100100001100110001110010101011";
                    when "00011" => level_vec_out <= "1011101111001001101011101110001101100100001100110001110010101011";
                    when "00100" => level_vec_out <= "1011101111001001101111101110001101100100001100110001110010111011";
                    when "00101" => level_vec_out <= "1011101111001001101111101110001101100100001100110101110010111011";
                    when "00110" => level_vec_out <= "1011101111001001101111101110001101100110001100110101110010111011";
                    when "00111" => level_vec_out <= "1011101111001001101111101110001101100110001100110101110010111011";
                    when "01000" => level_vec_out <= "1011101111001011101111101110001111100110011100110101110010111011";
                    when "01001" => level_vec_out <= "1011101111001011101111101110001111100110011110110111110010111011";
                    when "01010" => level_vec_out <= "1011101111001011101111101110101111100110011110110111110011111111";
                    when "01011" => level_vec_out <= "1011101111001011101111101110101111100110011110110111111011111111";
                    when "01100" => level_vec_out <= "1011101111001011101111101110101111100110011110110111111011111111";
                    when "01101" => level_vec_out <= "1011101111001011111111101110101111110111011110110111111011111111";
                    when "01110" => level_vec_out <= "1011101111001011111111101110101111111111011110110111111011111111";
                    when "01111" => level_vec_out <= "1011101111001011111111101110101111111111011110111111111011111111";
                    when "10000" => level_vec_out <= "1011111111101011111111101110101111111111011110111111111011111111";
                    when "10001" => level_vec_out <= "1011111111101011111111101110101111111111011110111111111011111111";
                    when "10010" => level_vec_out <= "1011111111101011111111101110101111111111011110111111111011111111";
                    when "10011" => level_vec_out <= "1011111111101011111111101110101111111111011110111111111011111111";
                    when "10100" => level_vec_out <= "1011111111101111111111101110101111111111011110111111111011111111";
                    when "10101" => level_vec_out <= "1011111111101111111111101110101111111111011110111111111011111111";
                    when "10110" => level_vec_out <= "1111111111101111111111101110101111111111011110111111111011111111";
                    when "10111" => level_vec_out <= "1111111111101111111111101110101111111111111110111111111011111111";
                    when "11000" => level_vec_out <= "1111111111101111111111101111101111111111111110111111111011111111";
                    when "11001" => level_vec_out <= "1111111111101111111111101111101111111111111110111111111011111111";
                    when "11010" => level_vec_out <= "1111111111101111111111101111101111111111111110111111111111111111";
                    when "11011" => level_vec_out <= "1111111111101111111111101111111111111111111110111111111111111111";
                    when "11100" => level_vec_out <= "1111111111101111111111101111111111111111111110111111111111111111";
                    when "11101" => level_vec_out <= "1111111111101111111111111111111111111111111111111111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "101" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1110100110001001101011100011110010101110001000110100001100110010";
                    when "00001" => level_vec_out <= "1110100110001001101111110011110010111110001100110100001100110010";
                    when "00010" => level_vec_out <= "1110100110001001101111110011110010111110001100110100001100110010";
                    when "00011" => level_vec_out <= "1110100110001101101111110011110010111110001100110100001100110010";
                    when "00100" => level_vec_out <= "1110100110001101101111110011110010111110001100110100001100110010";
                    when "00101" => level_vec_out <= "1110100110001101101111110011111010111110001100110100001100110010";
                    when "00110" => level_vec_out <= "1110100110001101101111110011111110111110001100110100001100110010";
                    when "00111" => level_vec_out <= "1111100110001101101111110011111110111110001100110110001110110110";
                    when "01000" => level_vec_out <= "1111100110001101101111110011111110111110001100110110001110110110";
                    when "01001" => level_vec_out <= "1111100110001101101111110011111110111110001100110110001110110110";
                    when "01010" => level_vec_out <= "1111100110001101101111110011111110111110001100110110001110110110";
                    when "01011" => level_vec_out <= "1111100110001101101111111011111110111110001100110110001110110110";
                    when "01100" => level_vec_out <= "1111100111001101101111111011111110111110001100110110001110110110";
                    when "01101" => level_vec_out <= "1111100111001101101111111011111110111110001100110110001110110110";
                    when "01110" => level_vec_out <= "1111100111001101101111111011111110111110011100110110001111110110";
                    when "01111" => level_vec_out <= "1111100111001101101111111011111110111110011100110110001111110110";
                    when "10000" => level_vec_out <= "1111100111001111101111111011111110111110011100110110001111110110";
                    when "10001" => level_vec_out <= "1111100111001111101111111011111111111110011100110110001111111110";
                    when "10010" => level_vec_out <= "1111100111001111101111111011111111111110011100110110101111111110";
                    when "10011" => level_vec_out <= "1111101111101111101111111011111111111110011100110110101111111110";
                    when "10100" => level_vec_out <= "1111101111101111101111111011111111111110011100110110101111111110";
                    when "10101" => level_vec_out <= "1111101111111111101111111011111111111110011101110111101111111110";
                    when "10110" => level_vec_out <= "1111101111111111111111111011111111111110011101110111101111111110";
                    when "10111" => level_vec_out <= "1111101111111111111111111011111111111110111101110111101111111110";
                    when "11000" => level_vec_out <= "1111101111111111111111111011111111111110111101110111101111111110";
                    when "11001" => level_vec_out <= "1111111111111111111111111011111111111110111111110111101111111110";
                    when "11010" => level_vec_out <= "1111111111111111111111111011111111111110111111111111101111111110";
                    when "11011" => level_vec_out <= "1111111111111111111111111011111111111111111111111111101111111110";
                    when "11100" => level_vec_out <= "1111111111111111111111111011111111111111111111111111101111111111";
                    when "11101" => level_vec_out <= "1111111111111111111111111011111111111111111111111111101111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111111111111111101111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "110" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0010100000111000100101111101010010011010011100100010100111110010";
                    when "00001" => level_vec_out <= "0010100001111000100101111101010010011010011100100010100111110010";
                    when "00010" => level_vec_out <= "0010101001111000100101111101010010011010011100100010100111110010";
                    when "00011" => level_vec_out <= "0010111001111000110101111101010010011010011100100011100111110011";
                    when "00100" => level_vec_out <= "0010111001111000110101111101010010011010011100100011100111110011";
                    when "00101" => level_vec_out <= "0010111001111100110101111111010010011010011100100011100111110011";
                    when "00110" => level_vec_out <= "1010111001111100110101111111010010011010011110100011110111110011";
                    when "00111" => level_vec_out <= "1010111001111100110101111111010010011110011110100011110111110011";
                    when "01000" => level_vec_out <= "1010111001111100110101111111010010011110011110100011110111110011";
                    when "01001" => level_vec_out <= "1010111001111100110101111111010010011110011110100011110111110011";
                    when "01010" => level_vec_out <= "1010111001111100110101111111010010011110011110100011110111110011";
                    when "01011" => level_vec_out <= "1010111001111100110101111111010010011110011110100011110111110011";
                    when "01100" => level_vec_out <= "1011111001111101110101111111010010111110011110100011110111110011";
                    when "01101" => level_vec_out <= "1011111001111111110101111111010010111110011110100011110111110011";
                    when "01110" => level_vec_out <= "1011111001111111110101111111011010111110111110100011110111110011";
                    when "01111" => level_vec_out <= "1011111001111111110101111111011010111110111110100011110111110011";
                    when "10000" => level_vec_out <= "1111111011111111110101111111011010111110111110100011110111110011";
                    when "10001" => level_vec_out <= "1111111011111111110101111111011010111110111110100011110111110011";
                    when "10010" => level_vec_out <= "1111111011111111110101111111011010111110111110101011110111110011";
                    when "10011" => level_vec_out <= "1111111011111111110101111111011010111110111110101011110111110011";
                    when "10100" => level_vec_out <= "1111111111111111110101111111011010111110111111101011110111110011";
                    when "10101" => level_vec_out <= "1111111111111111110101111111011010111110111111101011110111111011";
                    when "10110" => level_vec_out <= "1111111111111111110101111111011010111110111111101011111111111011";
                    when "10111" => level_vec_out <= "1111111111111111110101111111111011111111111111101011111111111111";
                    when "11000" => level_vec_out <= "1111111111111111110101111111111011111111111111101011111111111111";
                    when "11001" => level_vec_out <= "1111111111111111110101111111111011111111111111101011111111111111";
                    when "11010" => level_vec_out <= "1111111111111111110101111111111011111111111111101011111111111111";
                    when "11011" => level_vec_out <= "1111111111111111110111111111111011111111111111101011111111111111";
                    when "11100" => level_vec_out <= "1111111111111111111111111111111011111111111111101011111111111111";
                    when "11101" => level_vec_out <= "1111111111111111111111111111111011111111111111111011111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111011111111111111111011111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111011111111111111111011111111111111";
                when others => null;
                end case;
            when "111" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1010000011110010010001101000011111100111001000100101011000101110";
                    when "00001" => level_vec_out <= "1010000011110010010001101000011111100111001000100101011000101110";
                    when "00010" => level_vec_out <= "1010100011110010010001101000011111100111001000101101011000101110";
                    when "00011" => level_vec_out <= "1010100011110010010001101000011111100111001000101101011000111110";
                    when "00100" => level_vec_out <= "1010100011110010010001101000011111100111001000101101011000111110";
                    when "00101" => level_vec_out <= "1010100011110010010001101100011111100111001000101111011000111110";
                    when "00110" => level_vec_out <= "1010100111110010010001101100011111100111001000101111011000111110";
                    when "00111" => level_vec_out <= "1010100111110010010001101100011111100111001000101111011000111110";
                    when "01000" => level_vec_out <= "1011100111110010010001101100011111100111001100101111111000111110";
                    when "01001" => level_vec_out <= "1011100111110010010001101101011111100111001100101111111000111110";
                    when "01010" => level_vec_out <= "1011100111110010010001101101111111100111001100101111111010111110";
                    when "01011" => level_vec_out <= "1011100111110010010101101101111111100111001100101111111011111110";
                    when "01100" => level_vec_out <= "1011100111110010010101101101111111100111001100101111111011111110";
                    when "01101" => level_vec_out <= "1011100111110010010101101101111111100111001100101111111011111110";
                    when "01110" => level_vec_out <= "1011100111110010010101101101111111100111001100101111111011111110";
                    when "01111" => level_vec_out <= "1011100111110010011101101111111111110111001100101111111011111110";
                    when "10000" => level_vec_out <= "1011100111110010011101101111111111111111001100101111111011111110";
                    when "10001" => level_vec_out <= "1011100111110010011101101111111111111111001100101111111011111110";
                    when "10010" => level_vec_out <= "1011100111110010011111101111111111111111001100101111111011111110";
                    when "10011" => level_vec_out <= "1011100111110011011111101111111111111111001101101111111011111110";
                    when "10100" => level_vec_out <= "1011110111110011011111101111111111111111101101101111111011111110";
                    when "10101" => level_vec_out <= "1011110111110011111111101111111111111111101101101111111011111110";
                    when "10110" => level_vec_out <= "1011110111110011111111101111111111111111101101101111111011111110";
                    when "10111" => level_vec_out <= "1011110111110011111111101111111111111111101101101111111011111110";
                    when "11000" => level_vec_out <= "1111110111110011111111111111111111111111101101101111111011111110";
                    when "11001" => level_vec_out <= "1111110111110011111111111111111111111111101111111111111011111110";
                    when "11010" => level_vec_out <= "1111110111110011111111111111111111111111101111111111111111111110";
                    when "11011" => level_vec_out <= "1111110111110011111111111111111111111111101111111111111111111110";
                    when "11100" => level_vec_out <= "1111110111110011111111111111111111111111111111111111111111111110";
                    when "11101" => level_vec_out <= "1111110111110111111111111111111111111111111111111111111111111110";
                    when "11110" => level_vec_out <= "1111110111110111111111111111111111111111111111111111111111111110";
                    when "11111" => level_vec_out <= "1111110111110111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when others => null;
        end case;
    end process;
end Behavioral;