----
 -- @file level_hvec_gen_hdl.hpp
 -- @brief This script generates HDL code for generating high-dimensional LEVEL vectors.
 -- It is a novel method; for more information, please refer to our paper.
 --
 -- @author Saeid Jamili and Marco Angioli
 -- @note Author names are listed in alphabetical order.
 -- @email <saeid.jamili@uniroma1.it>
 -- @email <marco.angioli@uniroma1.it>
 --
 -- @contributors
 --
 -- @date Created: 24th July 2023
 -- @date Last Updated: 23th August 2023
 --
 -- @version 1.0.0
 --
 -- @institute Sapienza University of Rome
 -- @cite https://doi.org/10.xxxx/yyyyy
 --
 -- @section DEPENDENCIES
 -- - Dependency1: Description or version details.
 -- - Dependency2: Description or version details.
 --
 -- @section LICENSE
 -- This file is part of the Aeneas HyperCompute Platform.
 --
 -- Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 --
 -- @section CHANGELOG
 -- @version 1.0.0-dev - 23th August 2023
 -- - Initial release
 --
 -- @todo
 -- - Complete level vector generator function
 -- - Add training
 --
 -- @see
 -- -
 -- -
 -- -
 --
 --

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity level_vec_gen is
    Port ( level_vec_out : out  STD_LOGIC_VECTOR (63 downto 0);
           frame_index : in  STD_LOGIC_VECTOR (2 downto 0);
           frame_id : in  STD_LOGIC_VECTOR (4 downto 0));
end level_vec_gen;

architecture Behavioral of level_vec_gen is
begin
    process (frame_index, frame_id)
    begin
        -- Update this function to match your requirements
        case frame_index is
            when "000" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1000011101100110111100111000100101000001100010111000000101111110";
                    when "00001" => level_vec_out <= "1000011101100110111100111000100101010001100010111100000101111110";
                    when "00010" => level_vec_out <= "1000011101100110111100111000100101110001100010111100000101111110";
                    when "00011" => level_vec_out <= "1000011101100110111100111000100101110001100010111100000101111110";
                    when "00100" => level_vec_out <= "1010011101100110111100111000100101110001100010111100001101111110";
                    when "00101" => level_vec_out <= "1010011101100110111100111000100101110011100010111100001101111110";
                    when "00110" => level_vec_out <= "1010011101100110111100111000100101110011100010111100001101111110";
                    when "00111" => level_vec_out <= "1010011101100110111100111000100101110011100010111100001101111110";
                    when "01000" => level_vec_out <= "1110011101100110111100111000100101110011100010111100001101111110";
                    when "01001" => level_vec_out <= "1110011101100110111100111000110101110011100011111100001101111110";
                    when "01010" => level_vec_out <= "1110011101100110111100111000110111110011100011111100001101111110";
                    when "01011" => level_vec_out <= "1110011101100110111101111000110111110011100011111100001101111110";
                    when "01100" => level_vec_out <= "1110011101100110111101111000111111110011100011111100001101111110";
                    when "01101" => level_vec_out <= "1110011101100110111101111000111111110011100011111101001101111110";
                    when "01110" => level_vec_out <= "1110011101100110111101111000111111110011100011111101001101111110";
                    when "01111" => level_vec_out <= "1110011101100110111101111000111111110011100011111101101101111110";
                    when "10000" => level_vec_out <= "1110011101100110111101111001111111110011100011111101101101111110";
                    when "10001" => level_vec_out <= "1110011101100110111101111101111111110011100111111101101101111110";
                    when "10010" => level_vec_out <= "1110011111100110111101111101111111110011100111111101101111111110";
                    when "10011" => level_vec_out <= "1110111111100110111101111111111111110011100111111101101111111110";
                    when "10100" => level_vec_out <= "1110111111100110111101111111111111110011100111111101101111111110";
                    when "10101" => level_vec_out <= "1110111111100110111101111111111111110011100111111101101111111110";
                    when "10110" => level_vec_out <= "1110111111100110111111111111111111110011100111111101111111111110";
                    when "10111" => level_vec_out <= "1110111111100110111111111111111111110011100111111101111111111110";
                    when "11000" => level_vec_out <= "1110111111100110111111111111111111110011100111111101111111111110";
                    when "11001" => level_vec_out <= "1110111111100111111111111111111111110011100111111101111111111110";
                    when "11010" => level_vec_out <= "1110111111110111111111111111111111110011101111111101111111111110";
                    when "11011" => level_vec_out <= "1111111111110111111111111111111111110011101111111111111111111110";
                    when "11100" => level_vec_out <= "1111111111111111111111111111111111110011101111111111111111111110";
                    when "11101" => level_vec_out <= "1111111111111111111111111111111111111011111111111111111111111110";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111011111111111111111111111110";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "001" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1000111110011111011011001011000011111101111011101110101010110111";
                    when "00001" => level_vec_out <= "1000111110011111011011001011001011111101111011101110101010110111";
                    when "00010" => level_vec_out <= "1000111110011111011011001011001011111101111011111110101010110111";
                    when "00011" => level_vec_out <= "1000111110011111011011101011011111111101111011111110101010110111";
                    when "00100" => level_vec_out <= "1000111110011111011011101011011111111101111011111110101010110111";
                    when "00101" => level_vec_out <= "1000111110011111011011101011011111111101111011111111101010110111";
                    when "00110" => level_vec_out <= "1010111110011111011011101011011111111101111011111111101010110111";
                    when "00111" => level_vec_out <= "1011111110011111011011111011011111111101111011111111101010110111";
                    when "01000" => level_vec_out <= "1011111110011111011011111011011111111101111011111111101010110111";
                    when "01001" => level_vec_out <= "1011111110011111011011111011011111111101111011111111101010110111";
                    when "01010" => level_vec_out <= "1011111110011111011011111011011111111101111011111111101010110111";
                    when "01011" => level_vec_out <= "1011111110111111011011111011011111111101111011111111101010110111";
                    when "01100" => level_vec_out <= "1011111111111111011011111011011111111101111011111111101010110111";
                    when "01101" => level_vec_out <= "1111111111111111011011111011011111111101111011111111101010110111";
                    when "01110" => level_vec_out <= "1111111111111111011011111011011111111101111011111111101010110111";
                    when "01111" => level_vec_out <= "1111111111111111011011111011111111111101111011111111101010110111";
                    when "10000" => level_vec_out <= "1111111111111111011011111011111111111101111011111111101010110111";
                    when "10001" => level_vec_out <= "1111111111111111011011111011111111111101111011111111101010110111";
                    when "10010" => level_vec_out <= "1111111111111111011011111011111111111101111011111111101010110111";
                    when "10011" => level_vec_out <= "1111111111111111011011111011111111111101111011111111101010110111";
                    when "10100" => level_vec_out <= "1111111111111111011011111011111111111111111011111111101010110111";
                    when "10101" => level_vec_out <= "1111111111111111011011111011111111111111111011111111111010110111";
                    when "10110" => level_vec_out <= "1111111111111111011011111011111111111111111011111111111011110111";
                    when "10111" => level_vec_out <= "1111111111111111011011111011111111111111111011111111111011110111";
                    when "11000" => level_vec_out <= "1111111111111111011011111011111111111111111011111111111111110111";
                    when "11001" => level_vec_out <= "1111111111111111111111111011111111111111111011111111111111111111";
                    when "11010" => level_vec_out <= "1111111111111111111111111011111111111111111011111111111111111111";
                    when "11011" => level_vec_out <= "1111111111111111111111111011111111111111111011111111111111111111";
                    when "11100" => level_vec_out <= "1111111111111111111111111011111111111111111011111111111111111111";
                    when "11101" => level_vec_out <= "1111111111111111111111111011111111111111111011111111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111011111111111111111011111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111011111111111111111011111111111111111111";
                when others => null;
                end case;
            when "010" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1100000000001101011111111101111110001100100010110110011110010101";
                    when "00001" => level_vec_out <= "1100000000001111011111111101111110001100100010110110011110010101";
                    when "00010" => level_vec_out <= "1100000000001111011111111101111110001100100010110110011110010101";
                    when "00011" => level_vec_out <= "1100000000001111011111111101111110001110100010111110011110010101";
                    when "00100" => level_vec_out <= "1100000000001111011111111101111110001110100010111110011110010101";
                    when "00101" => level_vec_out <= "1100000000001111011111111101111110001110100010111110011110010101";
                    when "00110" => level_vec_out <= "1100000000001111011111111101111110001110100010111111111110010101";
                    when "00111" => level_vec_out <= "1100000000001111011111111101111110001110100010111111111110010101";
                    when "01000" => level_vec_out <= "1100100000001111011111111101111110001110100010111111111110110101";
                    when "01001" => level_vec_out <= "1100100000001111011111111101111110001110100010111111111110110101";
                    when "01010" => level_vec_out <= "1100100000001111011111111101111110001110100010111111111110110101";
                    when "01011" => level_vec_out <= "1100100000001111011111111101111110001110100010111111111110110101";
                    when "01100" => level_vec_out <= "1101100000001111011111111101111110001110100010111111111110110101";
                    when "01101" => level_vec_out <= "1101101000001111011111111101111110001110110010111111111110110101";
                    when "01110" => level_vec_out <= "1101101000001111011111111101111110001110110010111111111110110111";
                    when "01111" => level_vec_out <= "1101101000101111011111111101111110001110110010111111111110110111";
                    when "10000" => level_vec_out <= "1101101000101111011111111101111110001110110110111111111110110111";
                    when "10001" => level_vec_out <= "1101101000101111011111111101111110001110110110111111111110110111";
                    when "10010" => level_vec_out <= "1101101000101111011111111101111111001110110110111111111110110111";
                    when "10011" => level_vec_out <= "1101101010111111011111111101111111001110110110111111111110110111";
                    when "10100" => level_vec_out <= "1101101010111111011111111101111111001110110110111111111110110111";
                    when "10101" => level_vec_out <= "1101111010111111011111111101111111001110110110111111111110110111";
                    when "10110" => level_vec_out <= "1101111010111111011111111101111111001110110110111111111110111111";
                    when "10111" => level_vec_out <= "1101111110111111011111111101111111001110110110111111111110111111";
                    when "11000" => level_vec_out <= "1101111110111111011111111101111111001110110110111111111110111111";
                    when "11001" => level_vec_out <= "1101111110111111011111111101111111001110110110111111111110111111";
                    when "11010" => level_vec_out <= "1101111111111111011111111101111111011110110110111111111110111111";
                    when "11011" => level_vec_out <= "1111111111111111011111111101111111011110110110111111111110111111";
                    when "11100" => level_vec_out <= "1111111111111111111111111101111111011110110111111111111111111111";
                    when "11101" => level_vec_out <= "1111111111111111111111111101111111011111110111111111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111011111110111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111011111110111111111111111111111";
                when others => null;
                end case;
            when "011" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1000101000001111001000000001101011010100001110010010110000100111";
                    when "00001" => level_vec_out <= "1000101000001111001010000001101011110100001110010010110000100111";
                    when "00010" => level_vec_out <= "1000101000001111001010000001101011110100001110010010110000100111";
                    when "00011" => level_vec_out <= "1000101000001111001010000001101011110100001110010010110000100111";
                    when "00100" => level_vec_out <= "1100101010001111001010100001101011110100001110010010110000100111";
                    when "00101" => level_vec_out <= "1100101010001111001010100101101011110100001110010010110000100111";
                    when "00110" => level_vec_out <= "1100101010001111001010100101101011110100011110010010110000100111";
                    when "00111" => level_vec_out <= "1100101010001111101010100101101011110100011110010010111000100111";
                    when "01000" => level_vec_out <= "1100101010001111101010100101101011110100011110010010111000100111";
                    when "01001" => level_vec_out <= "1100101010001111101010100101101011110100011110010010111000100111";
                    when "01010" => level_vec_out <= "1100101010001111101010110101101011110100011110010010111100100111";
                    when "01011" => level_vec_out <= "1100101010001111101010110101101111110100011110010010111100100111";
                    when "01100" => level_vec_out <= "1100101010001111101010110101101111110100011110010010111100100111";
                    when "01101" => level_vec_out <= "1100101010001111101010110101101111110100011110010110111110100111";
                    when "01110" => level_vec_out <= "1100101010001111101011110101101111110100011110010110111110100111";
                    when "01111" => level_vec_out <= "1100101010001111101011110101101111110100011110010110111111100111";
                    when "10000" => level_vec_out <= "1100101010001111101011110101101111110100011110010110111111100111";
                    when "10001" => level_vec_out <= "1100101010001111101011111101101111110100011110010110111111100111";
                    when "10010" => level_vec_out <= "1100101010001111101011111101101111110110011110010110111111100111";
                    when "10011" => level_vec_out <= "1100101010001111101011111101101111110110011110010110111111100111";
                    when "10100" => level_vec_out <= "1110101010001111101111111101101111110110011110010110111111110111";
                    when "10101" => level_vec_out <= "1110101010001111101111111101101111110110011110110110111111111111";
                    when "10110" => level_vec_out <= "1110101010001111101111111101101111110110011110110110111111111111";
                    when "10111" => level_vec_out <= "1110101011001111101111111101101111110110011110110110111111111111";
                    when "11000" => level_vec_out <= "1110111011001111101111111101101111110110011111110110111111111111";
                    when "11001" => level_vec_out <= "1110111011001111101111111111101111110110011111110110111111111111";
                    when "11010" => level_vec_out <= "1110111011001111111111111111101111110110011111110110111111111111";
                    when "11011" => level_vec_out <= "1110111111101111111111111111101111110110011111110110111111111111";
                    when "11100" => level_vec_out <= "1110111111101111111111111111101111110111011111110110111111111111";
                    when "11101" => level_vec_out <= "1110111111101111111111111111101111110111011111110110111111111111";
                    when "11110" => level_vec_out <= "1111111111101111111111111111101111111111011111110111111111111111";
                    when "11111" => level_vec_out <= "1111111111101111111111111111111111111111011111110111111111111111";
                when others => null;
                end case;
            when "100" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1001010010000001000001110010000010010010100110001010001001001010";
                    when "00001" => level_vec_out <= "1001010010010001000001110010000010010010100110001010001001101010";
                    when "00010" => level_vec_out <= "1001010010010001100001110010000010010010100110001010001001111010";
                    when "00011" => level_vec_out <= "1001010010010001100001110010000010010010100110001010001001111010";
                    when "00100" => level_vec_out <= "1001010010010001100001110010000010010010100110001010001001111010";
                    when "00101" => level_vec_out <= "1001010010010101100001110010000010010010100111001110001001111010";
                    when "00110" => level_vec_out <= "1001010010010101100001110010000010010010100111001110001011111010";
                    when "00111" => level_vec_out <= "1001010010010101100001110010000010010010100111001110001011111010";
                    when "01000" => level_vec_out <= "1001010010010101100001110010000010110010100111011110001011111010";
                    when "01001" => level_vec_out <= "1001010010010101100101110010000010110010100111111110001011111010";
                    when "01010" => level_vec_out <= "1001011010010101100101110010000010110010100111111110001111111010";
                    when "01011" => level_vec_out <= "1001011010010101100111110010000010110011100111111110001111111010";
                    when "01100" => level_vec_out <= "1001011010010111100111110010010010110011100111111110101111111010";
                    when "01101" => level_vec_out <= "1001011010010111100111110010010010110011100111111110101111111010";
                    when "01110" => level_vec_out <= "1001011010110111100111110011010010110011100111111110101111111010";
                    when "01111" => level_vec_out <= "1001011011110111100111111011010010110011100111111110101111111010";
                    when "10000" => level_vec_out <= "1001011011110111100111111011010010110011100111111110101111111010";
                    when "10001" => level_vec_out <= "1001011011110111100111111011010010110011100111111110101111111010";
                    when "10010" => level_vec_out <= "1001011111110111100111111011010010110111100111111110101111111010";
                    when "10011" => level_vec_out <= "1001011111110111100111111011011010110111100111111110101111111110";
                    when "10100" => level_vec_out <= "1001011111110111100111111011111010110111100111111110101111111110";
                    when "10101" => level_vec_out <= "1001011111110111100111111011111010110111100111111110101111111110";
                    when "10110" => level_vec_out <= "1001011111110111101111111011111010110111100111111110101111111110";
                    when "10111" => level_vec_out <= "1001011111110111101111111111111010110111100111111110101111111110";
                    when "11000" => level_vec_out <= "1001011111110111111111111111111010111111100111111110101111111110";
                    when "11001" => level_vec_out <= "1001011111110111111111111111111011111111100111111110101111111111";
                    when "11010" => level_vec_out <= "1001011111110111111111111111111111111111100111111111101111111111";
                    when "11011" => level_vec_out <= "1001011111110111111111111111111111111111101111111111101111111111";
                    when "11100" => level_vec_out <= "1001011111110111111111111111111111111111111111111111101111111111";
                    when "11101" => level_vec_out <= "1011011111111111111111111111111111111111111111111111111111111111";
                    when "11110" => level_vec_out <= "1011111111111111111111111111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "101" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1110000000101001101100011010101111110001111010001101111000001001";
                    when "00001" => level_vec_out <= "1110000000101001101100011010101111110001111010001101111000001001";
                    when "00010" => level_vec_out <= "1110000000101001101101011010101111110001111010001101111000001001";
                    when "00011" => level_vec_out <= "1110000000101001101101011110101111110001111010001101111000001001";
                    when "00100" => level_vec_out <= "1110000000101001111101011110101111110001111010001101111000001001";
                    when "00101" => level_vec_out <= "1110000000101001111101011110101111110001111010001101111100001001";
                    when "00110" => level_vec_out <= "1110100000101001111101011110101111110001111010001101111100101001";
                    when "00111" => level_vec_out <= "1110100010101001111101011110101111110101111010001101111100101001";
                    when "01000" => level_vec_out <= "1110101010101001111101011110101111110111111110001101111100101001";
                    when "01001" => level_vec_out <= "1110101010101001111101011110101111110111111110011101111100101001";
                    when "01010" => level_vec_out <= "1110101010101001111101011110101111110111111110011111111100101001";
                    when "01011" => level_vec_out <= "1110101010101101111101011110101111111111111110011111111100101001";
                    when "01100" => level_vec_out <= "1110101010101101111101011110101111111111111110011111111100101001";
                    when "01101" => level_vec_out <= "1110101010101101111101011110101111111111111110011111111100101001";
                    when "01110" => level_vec_out <= "1110101010101101111101111110101111111111111110011111111100101001";
                    when "01111" => level_vec_out <= "1110101010101101111101111110101111111111111111011111111100101001";
                    when "10000" => level_vec_out <= "1110101011101101111111111110101111111111111111011111111100101001";
                    when "10001" => level_vec_out <= "1110101011101101111111111110101111111111111111011111111100101001";
                    when "10010" => level_vec_out <= "1110101011101101111111111110101111111111111111111111111100101001";
                    when "10011" => level_vec_out <= "1110101011101101111111111110101111111111111111111111111101101001";
                    when "10100" => level_vec_out <= "1110101011101111111111111110101111111111111111111111111101101001";
                    when "10101" => level_vec_out <= "1110101011101111111111111110101111111111111111111111111101101001";
                    when "10110" => level_vec_out <= "1110101011101111111111111110111111111111111111111111111101101001";
                    when "10111" => level_vec_out <= "1111101111101111111111111110111111111111111111111111111101101001";
                    when "11000" => level_vec_out <= "1111101111101111111111111111111111111111111111111111111101101001";
                    when "11001" => level_vec_out <= "1111101111101111111111111111111111111111111111111111111101101001";
                    when "11010" => level_vec_out <= "1111101111101111111111111111111111111111111111111111111101101101";
                    when "11011" => level_vec_out <= "1111101111101111111111111111111111111111111111111111111101101101";
                    when "11100" => level_vec_out <= "1111101111111111111111111111111111111111111111111111111111101101";
                    when "11101" => level_vec_out <= "1111101111111111111111111111111111111111111111111111111111101101";
                    when "11110" => level_vec_out <= "1111101111111111111111111111111111111111111111111111111111111101";
                    when "11111" => level_vec_out <= "1111101111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "110" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0000011101101100111101011001100000010111111100000101111100100110";
                    when "00001" => level_vec_out <= "0000011101101100111101011001100000010111111100000101111100100110";
                    when "00010" => level_vec_out <= "0001011101101100111101011001100000010111111100000101111100100110";
                    when "00011" => level_vec_out <= "0001011101101100111101011001100000110111111100000101111100100110";
                    when "00100" => level_vec_out <= "0001011101101100111101011011100000110111111100100101111100100110";
                    when "00101" => level_vec_out <= "0001011101101100111101011011100000110111111100100101111100100110";
                    when "00110" => level_vec_out <= "0001011101101100111101011011100000110111111100100101111100100110";
                    when "00111" => level_vec_out <= "1001011101101100111101011011100000110111111100100101111101100110";
                    when "01000" => level_vec_out <= "1001011101101100111101011011100000110111111100100101111101100110";
                    when "01001" => level_vec_out <= "1001011101101100111101011011100000110111111100100101111101110110";
                    when "01010" => level_vec_out <= "1001011101101101111101011011100000110111111100100101111101110110";
                    when "01011" => level_vec_out <= "1001011101101101111101011011110000110111111100100101111101110110";
                    when "01100" => level_vec_out <= "1001011101101101111101011011110001110111111100100101111101110110";
                    when "01101" => level_vec_out <= "1001011101101101111101011011110001110111111100100101111101111110";
                    when "01110" => level_vec_out <= "1001011101101101111101011011110001110111111100110101111101111110";
                    when "01111" => level_vec_out <= "1001011101101101111101011011110001110111111101110101111101111110";
                    when "10000" => level_vec_out <= "1001011101101111111101011011110001110111111101110101111101111110";
                    when "10001" => level_vec_out <= "1001111101101111111101011011110011110111111101110101111101111111";
                    when "10010" => level_vec_out <= "1001111101101111111101011011110011110111111101110101111101111111";
                    when "10011" => level_vec_out <= "1001111101101111111101011011110011110111111101111101111101111111";
                    when "10100" => level_vec_out <= "1001111101101111111101011011110011111111111101111101111101111111";
                    when "10101" => level_vec_out <= "1001111101111111111111011011110011111111111111111101111101111111";
                    when "10110" => level_vec_out <= "1001111111111111111111011011110011111111111111111101111101111111";
                    when "10111" => level_vec_out <= "1011111111111111111111011011110011111111111111111101111101111111";
                    when "11000" => level_vec_out <= "1011111111111111111111011011110011111111111111111111111111111111";
                    when "11001" => level_vec_out <= "1011111111111111111111011011110011111111111111111111111111111111";
                    when "11010" => level_vec_out <= "1011111111111111111111011011110011111111111111111111111111111111";
                    when "11011" => level_vec_out <= "1011111111111111111111011111110011111111111111111111111111111111";
                    when "11100" => level_vec_out <= "1011111111111111111111011111110011111111111111111111111111111111";
                    when "11101" => level_vec_out <= "1011111111111111111111011111111011111111111111111111111111111111";
                    when "11110" => level_vec_out <= "1011111111111111111111011111111011111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "111" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0000101111100111010111010011111000001011011001111110101010001110";
                    when "00001" => level_vec_out <= "0000101111100111010111010011111000001011011001111110101010001110";
                    when "00010" => level_vec_out <= "0000101111100111010111010011111000001111111001111110101010001110";
                    when "00011" => level_vec_out <= "0000101111100111010111010011111000001111111001111110101010101110";
                    when "00100" => level_vec_out <= "0000101111100111010111010011111000001111111001111110101010101110";
                    when "00101" => level_vec_out <= "0000101111100111010111010011111000001111111101111110101010101110";
                    when "00110" => level_vec_out <= "0000101111100111010111010011111000001111111101111110101011101110";
                    when "00111" => level_vec_out <= "0000101111100111010111010011111000001111111101111110101011101110";
                    when "01000" => level_vec_out <= "0000101111100111010111010011111000001111111101111110101011101110";
                    when "01001" => level_vec_out <= "0000101111100111010111010011111000001111111101111110101111101111";
                    when "01010" => level_vec_out <= "0000101111100111010111010011111000001111111101111110111111101111";
                    when "01011" => level_vec_out <= "0000101111100111010111010011111000001111111101111110111111101111";
                    when "01100" => level_vec_out <= "0001101111100111010111010011111000001111111101111110111111101111";
                    when "01101" => level_vec_out <= "1001101111100111010111010011111000001111111101111110111111101111";
                    when "01110" => level_vec_out <= "1001101111100111010111011111111000001111111101111110111111101111";
                    when "01111" => level_vec_out <= "1001101111100111010111011111111000001111111101111110111111101111";
                    when "10000" => level_vec_out <= "1001101111100111010111011111111011001111111101111111111111101111";
                    when "10001" => level_vec_out <= "1001101111111111010111011111111011001111111101111111111111101111";
                    when "10010" => level_vec_out <= "1001101111111111010111011111111011001111111111111111111111101111";
                    when "10011" => level_vec_out <= "1001101111111111010111011111111011001111111111111111111111101111";
                    when "10100" => level_vec_out <= "1101101111111111010111011111111011001111111111111111111111101111";
                    when "10101" => level_vec_out <= "1101101111111111010111011111111111001111111111111111111111101111";
                    when "10110" => level_vec_out <= "1101111111111111010111011111111111001111111111111111111111101111";
                    when "10111" => level_vec_out <= "1111111111111111110111011111111111001111111111111111111111101111";
                    when "11000" => level_vec_out <= "1111111111111111110111011111111111001111111111111111111111101111";
                    when "11001" => level_vec_out <= "1111111111111111110111011111111111101111111111111111111111101111";
                    when "11010" => level_vec_out <= "1111111111111111110111011111111111101111111111111111111111101111";
                    when "11011" => level_vec_out <= "1111111111111111111111011111111111101111111111111111111111101111";
                    when "11100" => level_vec_out <= "1111111111111111111111011111111111101111111111111111111111101111";
                    when "11101" => level_vec_out <= "1111111111111111111111111111111111101111111111111111111111101111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when others => null;
        end case;
    end process;
end Behavioral;