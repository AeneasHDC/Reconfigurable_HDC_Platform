----
 -- @file level_hvec_gen_hdl.hpp
 -- @brief This script generates HDL code for generating high-dimensional LEVEL vectors.
 -- It is a novel method; for more information, please refer to our paper.
 --
 -- @author Saeid Jamili and Marco Angioli
 -- @note Author names are listed in alphabetical order.
 -- @email <saeid.jamili@uniroma1.it>
 -- @email <marco.angioli@uniroma1.it>
 --
 -- @contributors
 --
 -- @date Created: 24th July 2023
 -- @date Last Updated: 23th August 2023
 --
 -- @version 0.0.1-dev
 --
 -- @institute Sapienza University of Rome
 -- @cite https://doi.org/10.xxxx/yyyyy
 --
 -- @section DEPENDENCIES
 -- - Dependency1: Description or version details.
 -- - Dependency2: Description or version details.
 --
 -- @section LICENSE
 -- This file is part of the Aeneas HyperCompute Platform.
 --
 -- Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 --
 -- @section CHANGELOG
 -- @version 1.0.0-dev - 23th August 2023
 -- - Initial release
 --
 -- @todo
 -- - Complete level vector generator function
 -- - Add training
 --
 -- @see
 -- -
 -- -
 -- -
 --
 --

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity level_vec_gen is
    Port ( level_vec_out : out  STD_LOGIC_VECTOR (99 downto 0);
           frame_index : in  STD_LOGIC_VECTOR (3 downto 0);
           frame_id : in  STD_LOGIC_VECTOR (4 downto 0));
end level_vec_gen;

architecture Behavioral of level_vec_gen is
begin
    process (frame_index, frame_id)
    begin
        -- Update this function to match your requirements
        case frame_index is
            when "0000" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0011100101100010100111001000010110101110010001010000100101110011010001011110011001010001100000111110";
                    when "00001" => level_vec_out <= "0011100101100010100111001000010110101110010001010000100101110011011001011110011011010001100000111110";
                    when "00010" => level_vec_out <= "0011100101100010100111001000010110101110010001010000100101110011011001011111011011011001100000111110";
                    when "00011" => level_vec_out <= "0011100101100010100111001000010110101110010001010000100101110011111001011111011011011001100000111110";
                    when "00100" => level_vec_out <= "0011100101100010100111001000010110101110010001010000100101110011111001011111011011011001100010111111";
                    when "00101" => level_vec_out <= "0011100101100010100111001100010110101110010001010000100101110011111001011111011011111001100010111111";
                    when "00110" => level_vec_out <= "0011110101100010100111001100010110101110010001010000100101110011111001011111011011111101100010111111";
                    when "00111" => level_vec_out <= "0011110101100010100111001100010110101110010001110000100101110011111001011111011011111101100010111111";
                    when "01000" => level_vec_out <= "0011110101100010100111001100010110101110110001110000100101110011111001011111011011111101100010111111";
                    when "01001" => level_vec_out <= "1011110101100010100111001100010110101110110001110000100101110011111001011111011011111101101010111111";
                    when "01010" => level_vec_out <= "1011110101100010100111001100010110101110110001110010100101110011111001011111011011111101101010111111";
                    when "01011" => level_vec_out <= "1011110101100010100111101100110110101110110011110010100101110011111001011111011011111101101010111111";
                    when "01100" => level_vec_out <= "1011110101100010100111101100110110101110110011110010100101110111111101011111011011111101101010111111";
                    when "01101" => level_vec_out <= "1011110101101010100111101100110110101110110011110010100101110111111101011111011111111101101011111111";
                    when "01110" => level_vec_out <= "1011110101101010101111101100110110101111110011110010100101110111111101011111011111111101101011111111";
                    when "01111" => level_vec_out <= "1011110101101010101111101100110110101111110011111010100101110111111101011111111111111101101011111111";
                    when "10000" => level_vec_out <= "1011110101111010101111101100110110101111110011111010100101111111111101011111111111111101101011111111";
                    when "10001" => level_vec_out <= "1011111101111010101111101100110110101111110011111010100101111111111101011111111111111101101011111111";
                    when "10010" => level_vec_out <= "1011111111111010101111101100110110101111110011111010110101111111111101011111111111111101101011111111";
                    when "10011" => level_vec_out <= "1011111111111010101111101100110110101111111011111010111101111111111111011111111111111101101011111111";
                    when "10100" => level_vec_out <= "1011111111111010101111101110110110101111111011111010111101111111111111011111111111111101101011111111";
                    when "10101" => level_vec_out <= "1011111111111010101111101110110110101111111011111010111101111111111111011111111111111101101011111111";
                    when "10110" => level_vec_out <= "1011111111111010101111101110110110101111111011111010111111111111111111011111111111111101101011111111";
                    when "10111" => level_vec_out <= "1011111111111010111111101110110110101111111111111010111111111111111111011111111111111101101011111111";
                    when "11000" => level_vec_out <= "1011111111111010111111101110111110101111111111111010111111111111111111011111111111111101101111111111";
                    when "11001" => level_vec_out <= "1011111111111110111111101110111110101111111111111010111111111111111111111111111111111101101111111111";
                    when "11010" => level_vec_out <= "1011111111111110111111101110111110101111111111111011111111111111111111111111111111111101101111111111";
                    when "11011" => level_vec_out <= "1011111111111110111111101110111111101111111111111011111111111111111111111111111111111101111111111111";
                    when "11100" => level_vec_out <= "1111111111111110111111101110111111101111111111111111111111111111111111111111111111111111111111111111";
                    when "11101" => level_vec_out <= "1111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "0001" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1000011000010101010110001011010100010000100101100110111110001101111100101110101111001110011111101100";
                    when "00001" => level_vec_out <= "1100011001010101010110001011010100010000100101100110111110001101111100101110101111001110011111101100";
                    when "00010" => level_vec_out <= "1100011001010101010110101011010100010000100111100110111110001101111100101110101111001110011111101100";
                    when "00011" => level_vec_out <= "1100011001010101010110101011010100010000100111100110111110001101111100101110101111011111011111101100";
                    when "00100" => level_vec_out <= "1101011001010101010110101011010100010000100111100110111110101101111100101110101111011111011111101100";
                    when "00101" => level_vec_out <= "1101111001010101010110101011011100010000100111100110111110101101111100101110101111011111011111101100";
                    when "00110" => level_vec_out <= "1101111001010101010110101011011100010000100111100110111110101101111100101110101111011111011111101100";
                    when "00111" => level_vec_out <= "1101111001010101010111101011011100010000100111100110111110101101111100101110101111011111011111101100";
                    when "01000" => level_vec_out <= "1101111001010101010111101011011100010000100111100110111110101101111100101110101111011111111111101100";
                    when "01001" => level_vec_out <= "1101111011010101010111101011011100010000100111100110111110101101111100101110101111011111111111101100";
                    when "01010" => level_vec_out <= "1101111011010101010111101011011100010000100111100110111110101101111100101110101111011111111111101100";
                    when "01011" => level_vec_out <= "1101111011010101010111101011011100010000100111100110111110101101111100101110101111011111111111101100";
                    when "01100" => level_vec_out <= "1101111011010101010111101011011100010010100111100110111110101101111100101110101111011111111111101100";
                    when "01101" => level_vec_out <= "1101111011010101010111101011011100010010100111100110111110101101111100101110101111011111111111101100";
                    when "01110" => level_vec_out <= "1101111011011101010111101011011100010010100111100110111110101101111100101110101111111111111111101100";
                    when "01111" => level_vec_out <= "1101111011011101010111101011011100010010100111100110111110101101111100101110101111111111111111101100";
                    when "10000" => level_vec_out <= "1101111011011101010111101011011110010110100111100110111110101101111100101110101111111111111111101100";
                    when "10001" => level_vec_out <= "1101111011011101010111101011011110011110100111100110111110101101111100101110101111111111111111101100";
                    when "10010" => level_vec_out <= "1101111011011101011111101011011110011110100111100110111110101101111100101110101111111111111111101100";
                    when "10011" => level_vec_out <= "1101111011011101011111101011011110011110100111100110111111101101111100101110101111111111111111101100";
                    when "10100" => level_vec_out <= "1101111011011101011111101011111110011110100111100110111111101101111100101110101111111111111111101110";
                    when "10101" => level_vec_out <= "1101111011011101111111101011111110011110100111100110111111101101111100101110101111111111111111101110";
                    when "10110" => level_vec_out <= "1101111111111101111111101011111110011110100111100110111111101101111100101110101111111111111111101110";
                    when "10111" => level_vec_out <= "1101111111111111111111101111111110011110100111100111111111101101111110101110101111111111111111101110";
                    when "11000" => level_vec_out <= "1101111111111111111111101111111110011111100111100111111111101101111110101111101111111111111111101110";
                    when "11001" => level_vec_out <= "1111111111111111111111101111111110011111101111100111111111101101111110111111101111111111111111101111";
                    when "11010" => level_vec_out <= "1111111111111111111111101111111110011111101111110111111111101101111110111111101111111111111111101111";
                    when "11011" => level_vec_out <= "1111111111111111111111111111111110111111101111110111111111101101111110111111101111111111111111101111";
                    when "11100" => level_vec_out <= "1111111111111111111111111111111110111111101111110111111111101101111110111111101111111111111111111111";
                    when "11101" => level_vec_out <= "1111111111111111111111111111111111111111101111110111111111101101111111111111101111111111111111111111";
                when others => null;
                end case;
            when "0010" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0100010100011101001000010001100111011001000110010111011000100010100111110111100110011001100111100011";
                    when "00001" => level_vec_out <= "0100010100011101001000010011100111011001000110010111011000100010100111110111100110011001100111100011";
                    when "00010" => level_vec_out <= "0100010100011101001000010011100111011001000110010111011100100010100111110111100110011001100111100011";
                    when "00011" => level_vec_out <= "0100010100011101001000010011100111011001000110010111011100100010100111110111100110011001100111100011";
                    when "00100" => level_vec_out <= "0100010100011101001000010011100111011001000110010111011100100010100111110111100110011001100111100011";
                    when "00101" => level_vec_out <= "0100010100011101001000010011100111011001000110110111011100100010100111110111100110011001100111101011";
                    when "00110" => level_vec_out <= "0100010110011101001000010011100111011001000111110111011100100010100111110111100110011101100111101011";
                    when "00111" => level_vec_out <= "0100010110011101001000110011100111011001000111110111011100100010100111110111100110011101100111101011";
                    when "01000" => level_vec_out <= "0100010110011101001000110011100111011001000111110111011100100010100111110111100110011101100111101011";
                    when "01001" => level_vec_out <= "0100010110011101001000110011100111011001000111110111011100100010100111110111100110011101100111101011";
                    when "01010" => level_vec_out <= "0100010110011101101000110011100111011001000111110111011100101010100111110111100110011101100111101011";
                    when "01011" => level_vec_out <= "0100110110011101101000110011110111011001000111110111011100101010100111110111100110011101100111101011";
                    when "01100" => level_vec_out <= "0100110110011101101000110011110111011001001111110111011100101010110111110111100111011101100111101111";
                    when "01101" => level_vec_out <= "0100110110011101101000110011110111011001001111110111011100101010110111110111100111011101100111101111";
                    when "01110" => level_vec_out <= "0100110110011101101000110011110111011001001111110111111100101010110111110111100111011101100111101111";
                    when "01111" => level_vec_out <= "0100110110011101101000110011110111011001001111110111111100101010110111110111100111011101100111101111";
                    when "10000" => level_vec_out <= "0100110110011101101000110011110111011001001111110111111100101010110111110111100111011101100111101111";
                    when "10001" => level_vec_out <= "0100110110011101101000110011110111111001001111110111111100101010110111110111110111011101100111101111";
                    when "10010" => level_vec_out <= "0101110110011101101000110011110111111001001111111111111110101110110111110111110111011111100111101111";
                    when "10011" => level_vec_out <= "1101111110011101101000110011111111111011001111111111111110101110110111110111111111011111100111101111";
                    when "10100" => level_vec_out <= "1101111110011101101000110011111111111011001111111111111110111110110111111111111111111111100111101111";
                    when "10101" => level_vec_out <= "1101111110011101101000110011111111111011001111111111111110111110111111111111111111111111100111101111";
                    when "10110" => level_vec_out <= "1101111110011101101000110011111111111011001111111111111110111110111111111111111111111111100111101111";
                    when "10111" => level_vec_out <= "1101111110011111101000110011111111111111001111111111111110111110111111111111111111111111100111101111";
                    when "11000" => level_vec_out <= "1101111110011111101000110011111111111111101111111111111110111110111111111111111111111111100111101111";
                    when "11001" => level_vec_out <= "1101111110011111101000110011111111111111111111111111111110111110111111111111111111111111101111101111";
                    when "11010" => level_vec_out <= "1101111110011111101101110011111111111111111111111111111111111110111111111111111111111111111111101111";
                    when "11011" => level_vec_out <= "1101111110011111101101111011111111111111111111111111111111111111111111111111111111111111111111101111";
                    when "11100" => level_vec_out <= "1101111110011111101101111011111111111111111111111111111111111111111111111111111111111111111111101111";
                    when "11101" => level_vec_out <= "1111111111011111101101111011111111111111111111111111111111111111111111111111111111111111111111101111";
                when others => null;
                end case;
            when "0011" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1110100001011101100011001010011101101000100111100100010101101011111001101001111001101100010111100010";
                    when "00001" => level_vec_out <= "1110100001011101100011001010011101101000100111100100010101101011111001101001111001101100010111100010";
                    when "00010" => level_vec_out <= "1110100001011101100011001010011101101000100111100100010101101011111001101001111001101100010111100010";
                    when "00011" => level_vec_out <= "1110100001011101100011001010011101101000100111100100010101101011111001101001111001101101010111100110";
                    when "00100" => level_vec_out <= "1111101001011101100011001010011101101010100111100100010101101011111001101001111001101101010111100111";
                    when "00101" => level_vec_out <= "1111101001011101100011001010011101101010100111100100010101101011111001101001111001101101010111101111";
                    when "00110" => level_vec_out <= "1111101001111101100011001010011101101010100111100101010101101011111001101001111001101101011111101111";
                    when "00111" => level_vec_out <= "1111101001111101101011001010011101101010100111100101010101101011111001101101111001101101011111101111";
                    when "01000" => level_vec_out <= "1111111001111101101011001010011101101010100111100101010101101011111001101101111001101101011111101111";
                    when "01001" => level_vec_out <= "1111111001111101101011001010111101101010100111100101010101101011111011101101111001101101011111101111";
                    when "01010" => level_vec_out <= "1111111001111101101011001010111101101011100111100101010101101011111011101101111001101101011111101111";
                    when "01011" => level_vec_out <= "1111111001111101101011001010111101101011100111100101010101101011111011101111111001101101011111101111";
                    when "01100" => level_vec_out <= "1111111001111101101011001010111101101011100111100101010101101011111011101111111001101101011111101111";
                    when "01101" => level_vec_out <= "1111111001111101101011001010111101111011100111100101010101101011111011101111111001101111011111101111";
                    when "01110" => level_vec_out <= "1111111001111101101011001010111101111011100111110101010101101011111011101111111001101111111111101111";
                    when "01111" => level_vec_out <= "1111111001111101111011001010111101111011100111110101010111101111111011101111111001111111111111101111";
                    when "10000" => level_vec_out <= "1111111011111101111011111010111101111111100111110101010111101111111011101111111011111111111111111111";
                    when "10001" => level_vec_out <= "1111111011111111111011111010111101111111110111110101010111101111111011101111111011111111111111111111";
                    when "10010" => level_vec_out <= "1111111011111111111011111010111101111111110111110101010111101111111011111111111111111111111111111111";
                    when "10011" => level_vec_out <= "1111111011111111111011111010111101111111110111110101010111101111111011111111111111111111111111111111";
                    when "10100" => level_vec_out <= "1111111011111111111011111011111101111111111111110101010111101111111011111111111111111111111111111111";
                    when "10101" => level_vec_out <= "1111111011111111111011111011111101111111111111110101010111101111111011111111111111111111111111111111";
                    when "10110" => level_vec_out <= "1111111011111111111011111011111101111111111111110101010111101111111011111111111111111111111111111111";
                    when "10111" => level_vec_out <= "1111111011111111111011111011111101111111111111110101110111101111111011111111111111111111111111111111";
                    when "11000" => level_vec_out <= "1111111011111111111011111111111101111111111111110101110111101111111011111111111111111111111111111111";
                    when "11001" => level_vec_out <= "1111111011111111111011111111111101111111111111110101111111111111111011111111111111111111111111111111";
                    when "11010" => level_vec_out <= "1111111011111111111011111111111101111111111111110111111111111111111011111111111111111111111111111111";
                    when "11011" => level_vec_out <= "1111111111111111111111111111111101111111111111110111111111111111111011111111111111111111111111111111";
                    when "11100" => level_vec_out <= "1111111111111111111111111111111111111111111111110111111111111111111011111111111111111111111111111111";
                    when "11101" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111";
                when others => null;
                end case;
            when "0100" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0100000110110111001011000001101001001101110001001101011111001110000011011111000110110001011010011111";
                    when "00001" => level_vec_out <= "0100000110110111001011000001101001001101110001001101011111001110000011011111000110110001011111011111";
                    when "00010" => level_vec_out <= "0100000110110111001011000001101101001101110001001101011111001110000011011111000110110001011111011111";
                    when "00011" => level_vec_out <= "0100000110110111101011000001101101001101110001001101011111001110000011011111000110110001011111011111";
                    when "00100" => level_vec_out <= "0100000110110111101011000101101101001101110001001101011111001110000011011111000110110001011111011111";
                    when "00101" => level_vec_out <= "0100000110110111101011000101101101001101110001001101011111001110000011011111000110110001011111011111";
                    when "00110" => level_vec_out <= "0100000110110111101011000101101101001101110001001101011111101110000011011111001110110001011111011111";
                    when "00111" => level_vec_out <= "0100010110110111101011000101101101001101110001001111011111101110000011011111001110110001011111011111";
                    when "01000" => level_vec_out <= "1100010110110111101011000101101101001101110001001111111111101110100011011111001110110001011111111111";
                    when "01001" => level_vec_out <= "1100010110110111101011000101101101001101110001001111111111101110100011011111001110110001011111111111";
                    when "01010" => level_vec_out <= "1100010110110111101011000101101101001101110001001111111111101110101011011111001110110001011111111111";
                    when "01011" => level_vec_out <= "1100010110110111101011000101101101001101110001001111111111101110101011011111001110110001011111111111";
                    when "01100" => level_vec_out <= "1100010110110111101011000101101101001101110001001111111111101110101011011111101110110001011111111111";
                    when "01101" => level_vec_out <= "1100010110110111101011000101101101001101110001001111111111101110101011011111101110110001011111111111";
                    when "01110" => level_vec_out <= "1100110110110111101011000101101101011101110001001111111111101110101011011111101110110101011111111111";
                    when "01111" => level_vec_out <= "1100110110110111101011000101101101011101110001101111111111101110101011011111101110110101011111111111";
                    when "10000" => level_vec_out <= "1101110110110111101011000101101101011101110001101111111111101110101011011111101110110101011111111111";
                    when "10001" => level_vec_out <= "1101110110110111101111000101101101011101110001101111111111101111101011011111101111110101011111111111";
                    when "10010" => level_vec_out <= "1101110110110111101111000101101101011101110001101111111111101111101011011111101111110101011111111111";
                    when "10011" => level_vec_out <= "1101110110111111101111000101101101011101110001101111111111101111101011011111101111110101011111111111";
                    when "10100" => level_vec_out <= "1111110110111111101111000101101101011101111001101111111111101111111011011111101111110101011111111111";
                    when "10101" => level_vec_out <= "1111110110111111101111100101111101011101111101101111111111101111111011011111101111111101011111111111";
                    when "10110" => level_vec_out <= "1111111110111111101111100101111101011101111101101111111111111111111011011111101111111101111111111111";
                    when "10111" => level_vec_out <= "1111111110111111101111110101111101011101111101111111111111111111111011011111101111111101111111111111";
                    when "11000" => level_vec_out <= "1111111110111111101111110111111101011111111101111111111111111111111011011111101111111101111111111111";
                    when "11001" => level_vec_out <= "1111111110111111101111110111111101011111111101111111111111111111111011011111101111111111111111111111";
                    when "11010" => level_vec_out <= "1111111110111111111111110111111101011111111101111111111111111111111011011111111111111111111111111111";
                    when "11011" => level_vec_out <= "1111111110111111111111110111111101111111111101111111111111111111111011011111111111111111111111111111";
                    when "11100" => level_vec_out <= "1111111110111111111111110111111101111111111101111111111111111111111011011111111111111111111111111111";
                    when "11101" => level_vec_out <= "1111111110111111111111110111111101111111111101111111111111111111111011011111111111111111111111111111";
                when others => null;
                end case;
            when "0101" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1010110000010000110100010000101110010100010010000000001110011100001101011010000000000000010000001000";
                    when "00001" => level_vec_out <= "1010110000010000110100010000101110010100010010000000001110011101001101011010000000000100010001001000";
                    when "00010" => level_vec_out <= "1010110000010000111100110000101110010100010010000000011110011101001111011010000000100100010001001000";
                    when "00011" => level_vec_out <= "1010110000010000111100110000101110010100010010000000011110011101001111011010000000100100010001001000";
                    when "00100" => level_vec_out <= "1010110000010000111100110000101110010110010010000000011110011101001111011010100000100100010001001000";
                    when "00101" => level_vec_out <= "1010110000010000111100110000101110010110010010000000111110011101001111011010100000100101010011001000";
                    when "00110" => level_vec_out <= "1010110000010000111100110001101110010110010010010000111110011101001111011010100000100101010011001000";
                    when "00111" => level_vec_out <= "1010110000010000111100110001101110010110010110110000111110011101001111011010100000100101010011001100";
                    when "01000" => level_vec_out <= "1010110000010000111100110001101110010110010111110000111110011101001111011010110100100101010011001101";
                    when "01001" => level_vec_out <= "1010110001110000111101110001101110010110010111110000111110011101001111011010110101100101110011001101";
                    when "01010" => level_vec_out <= "1010110101110001111111110001101110010110010111110000111110011101001111011010110101100101110011001101";
                    when "01011" => level_vec_out <= "1010110111110001111111110001101110010110010111110000111111011101101111011010110101110101110011001101";
                    when "01100" => level_vec_out <= "1010110111110001111111110001101110010110010111110000111111011101101111011010110101110101110111001101";
                    when "01101" => level_vec_out <= "1010110111110001111111110001101110010110010111110000111111011101101111011010111101110111110111001101";
                    when "01110" => level_vec_out <= "1010110111110101111111110001101110110110010111110000111111011101101111011010111101110111110111001101";
                    when "01111" => level_vec_out <= "1010110111110101111111110001101110110110011111110000111111011101101111011010111101110111110111001101";
                    when "10000" => level_vec_out <= "1010110111110101111111110001101110110110011111110000111111011101101111011010111101110111110111001101";
                    when "10001" => level_vec_out <= "1010110111110101111111110001101110110111011111110000111111011101101111011010111101110111110111001101";
                    when "10010" => level_vec_out <= "1010110111111101111111111001101110110111011111110000111111011101101111011010111101110111110111001101";
                    when "10011" => level_vec_out <= "1010110111111111111111111001101110110111011111110000111111011101101111011110111101110111110111001101";
                    when "10100" => level_vec_out <= "1010110111111111111111111001101110110111011111110001111111011101101111011111111101110111110111001101";
                    when "10101" => level_vec_out <= "1011110111111111111111111001101110110111011111110001111111011101101111011111111101110111110111101101";
                    when "10110" => level_vec_out <= "1111110111111111111111111101101110110111011111110001111111011101101111111111111101110111110111101111";
                    when "10111" => level_vec_out <= "1111110111111111111111111101101110110111011111110001111111011101101111111111111101110111110111101111";
                    when "11000" => level_vec_out <= "1111110111111111111111111101101110110111011111110001111111111101101111111111111111111111110111101111";
                    when "11001" => level_vec_out <= "1111110111111111111111111101111110110111011111110001111111111101101111111111111111111111110111101111";
                    when "11010" => level_vec_out <= "1111110111111111111111111111111110110111011111110001111111111101101111111111111111111111110111101111";
                    when "11011" => level_vec_out <= "1111110111111111111111111111111110110111011111110001111111111101101111111111111111111111110111101111";
                    when "11100" => level_vec_out <= "1111110111111111111111111111111111111111111111110001111111111101101111111111111111111111110111101111";
                    when "11101" => level_vec_out <= "1111110111111111111111111111111111111111111111110101111111111101101111111111111111111111111111101111";
                when others => null;
                end case;
            when "0110" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1110101011000011110010111111010110110111111111111101000101111100100100100011010011101111111000011111";
                    when "00001" => level_vec_out <= "1110111011000011110010111111010110110111111111111101000101111100100100100011010011101111111000011111";
                    when "00010" => level_vec_out <= "1110111011000111110010111111010110110111111111111101000101111100100100100011010011101111111000011111";
                    when "00011" => level_vec_out <= "1110111011100111110010111111010110110111111111111101010101111100100100100011010011101111111000011111";
                    when "00100" => level_vec_out <= "1110111011100111110010111111010110110111111111111101010101111100100100100011010011101111111000011111";
                    when "00101" => level_vec_out <= "1110111011100111110010111111010110110111111111111101010101111100100101100011011011101111111000011111";
                    when "00110" => level_vec_out <= "1110111011101111110010111111010110110111111111111101010101111100100101101011011011101111111000011111";
                    when "00111" => level_vec_out <= "1110111011101111110110111111010110110111111111111101010101111101100101101011011011101111111000011111";
                    when "01000" => level_vec_out <= "1110111011101111110110111111010110110111111111111101010101111101101101101011011011101111111000011111";
                    when "01001" => level_vec_out <= "1110111011101111110110111111010110110111111111111101010101111101101101101011011011111111111000011111";
                    when "01010" => level_vec_out <= "1110111011101111110110111111010110110111111111111101010101111101101101101011011011111111111001011111";
                    when "01011" => level_vec_out <= "1110111011101111110110111111010110110111111111111101010101111101101101111011011011111111111001011111";
                    when "01100" => level_vec_out <= "1110111011101111110110111111010110110111111111111101010101111111101101111011011011111111111001011111";
                    when "01101" => level_vec_out <= "1110111111111111110110111111010110110111111111111101010101111111101101111011011011111111111001011111";
                    when "01110" => level_vec_out <= "1110111111111111110110111111010110110111111111111101010101111111101111111011011011111111111001011111";
                    when "01111" => level_vec_out <= "1110111111111111110110111111010110110111111111111101010101111111101111111011011011111111111001111111";
                    when "10000" => level_vec_out <= "1110111111111111110110111111010110110111111111111101010101111111101111111011011011111111111001111111";
                    when "10001" => level_vec_out <= "1110111111111111110110111111010110110111111111111101010101111111101111111011011011111111111001111111";
                    when "10010" => level_vec_out <= "1110111111111111110110111111010110110111111111111101110101111111101111111011011011111111111001111111";
                    when "10011" => level_vec_out <= "1110111111111111110110111111010110110111111111111101110101111111101111111011011011111111111001111111";
                    when "10100" => level_vec_out <= "1110111111111111110110111111010110110111111111111101110101111111101111111011011011111111111001111111";
                    when "10101" => level_vec_out <= "1110111111111111110110111111010110110111111111111101110101111111101111111011011011111111111011111111";
                    when "10110" => level_vec_out <= "1110111111111111110111111111010110110111111111111101110101111111111111111111011111111111111011111111";
                    when "10111" => level_vec_out <= "1110111111111111110111111111010110110111111111111101110111111111111111111111011111111111111011111111";
                    when "11000" => level_vec_out <= "1110111111111111111111111111010110110111111111111101110111111111111111111111011111111111111011111111";
                    when "11001" => level_vec_out <= "1110111111111111111111111111010110111111111111111101110111111111111111111111011111111111111011111111";
                    when "11010" => level_vec_out <= "1110111111111111111111111111010110111111111111111101110111111111111111111111011111111111111111111111";
                    when "11011" => level_vec_out <= "1110111111111111111111111111010110111111111111111101111111111111111111111111011111111111111111111111";
                    when "11100" => level_vec_out <= "1111111111111111111111111111010110111111111111111111111111111111111111111111111111111111111111111111";
                    when "11101" => level_vec_out <= "1111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "0111" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0001111000101111110100011111100001000110011000010101100111100101100111010101011001011100001001111101";
                    when "00001" => level_vec_out <= "0101111000101111110100011111100001000110011000010101100111100101100111010101011001011100001001111111";
                    when "00010" => level_vec_out <= "0101111000101111110100011111100111000110011000010101100111100101100111010101011001011100001001111111";
                    when "00011" => level_vec_out <= "0101111000101111110100011111100111000110011000010101100111100101100111010101111001011100001001111111";
                    when "00100" => level_vec_out <= "0101111000101111110100011111100111000110011000010101100111100101100111010101111001011100001001111111";
                    when "00101" => level_vec_out <= "0111111000101111110100011111100111000110011000010101100111100101110111010101111001011100001001111111";
                    when "00110" => level_vec_out <= "0111111000101111110100011111100111000110011000010101100111100101110111010101111001011100001001111111";
                    when "00111" => level_vec_out <= "0111111000101111110100011111100111100110011000010101100111100101110111010101111101011100001001111111";
                    when "01000" => level_vec_out <= "0111111001101111110100011111100111100110011000010101100111100101110111010101111101011100001001111111";
                    when "01001" => level_vec_out <= "0111111001101111110100011111100111110110011000010101100111100101110111010101111101011100001001111111";
                    when "01010" => level_vec_out <= "0111111001101111110100011111100111110110011000010101100111100101110111010101111101011100101001111111";
                    when "01011" => level_vec_out <= "0111111001101111110100011111100111111110011010110101100111110101110111010101111101011100101001111111";
                    when "01100" => level_vec_out <= "0111111001101111110100011111100111111110011010111101100111110101110111010101111101011100101001111111";
                    when "01101" => level_vec_out <= "0111111001101111110100011111100111111110011010111101100111111101110111010101111101011101101001111111";
                    when "01110" => level_vec_out <= "0111111001101111110100011111100111111110011010111101100111111101110111010101111101011101101011111111";
                    when "01111" => level_vec_out <= "0111111001101111110100011111100111111110011010111101100111111101111111010101111101011101101011111111";
                    when "10000" => level_vec_out <= "0111111001101111110100011111100111111110011011111101100111111101111111110101111101011101101011111111";
                    when "10001" => level_vec_out <= "0111111001101111110100111111100111111110011011111101100111111101111111111101111101011101101011111111";
                    when "10010" => level_vec_out <= "0111111001101111110100111111100111111110011011111101100111111101111111111101111101011101101011111111";
                    when "10011" => level_vec_out <= "0111111001101111110101111111100111111110011011111101100111111101111111111111111101011101101011111111";
                    when "10100" => level_vec_out <= "0111111001101111110111111111100111111110011011111101100111111101111111111111111101011101101011111111";
                    when "10101" => level_vec_out <= "1111111001101111110111111111100111111110011011111101100111111101111111111111111101011101101011111111";
                    when "10110" => level_vec_out <= "1111111001101111110111111111100111111110011011111101100111111101111111111111111101011101101011111111";
                    when "10111" => level_vec_out <= "1111111001101111110111111111100111111110111011111101100111111101111111111111111101011101101011111111";
                    when "11000" => level_vec_out <= "1111111001101111110111111111100111111111111111111101100111111101111111111111111101011101101011111111";
                    when "11001" => level_vec_out <= "1111111001111111110111111111100111111111111111111101100111111101111111111111111101011111101011111111";
                    when "11010" => level_vec_out <= "1111111101111111110111111111100111111111111111111101100111111101111111111111111101111111101011111111";
                    when "11011" => level_vec_out <= "1111111101111111110111111111101111111111111111111101101111111101111111111111111101111111101011111111";
                    when "11100" => level_vec_out <= "1111111101111111111111111111111111111111111111111111111111111101111111111111111101111111111011111111";
                    when "11101" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111011111111";
                when others => null;
                end case;
            when "1000" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0011110000111111001000001111100011100011110010110101000010001111110010000110100001101011100001010000";
                    when "00001" => level_vec_out <= "0011110000111111001000011111100011100011110010110101000010001111110010000110100001101011100001010000";
                    when "00010" => level_vec_out <= "0011110000111111001000011111100011100011110010110101000010001111110010000110100001101011100001010000";
                    when "00011" => level_vec_out <= "0011110000111111001000011111101111100011110010110101001010001111110010000110100001101011100001010000";
                    when "00100" => level_vec_out <= "1011110000111111001000011111101111100011110010110101001010001111110010000110100001101011100001010101";
                    when "00101" => level_vec_out <= "1011110000111111001000011111101111100011110010110101001010001111110010000110100001101011100001010101";
                    when "00110" => level_vec_out <= "1011110000111111001000011111101111100011111010110101001010001111110010000110100001101011100001010101";
                    when "00111" => level_vec_out <= "1011110000111111001000011111101111100011111010111101001010001111110010000110100001101011100001010101";
                    when "01000" => level_vec_out <= "1011110000111111001000011111101111100011111010111101001010001111110010000110100001101011101101010101";
                    when "01001" => level_vec_out <= "1011110000111111001100011111101111100011111010111101001010011111110110000110100001101011101101010101";
                    when "01010" => level_vec_out <= "1011110001111111001100011111101111100011111011111101001110011111110110000110111001101011101101110101";
                    when "01011" => level_vec_out <= "1011110001111111001100011111101111100011111011111101001110011111110110000110111001101011101101110101";
                    when "01100" => level_vec_out <= "1011110001111111001100011111101111100011111011111101001110011111110110001110111001111011111101110101";
                    when "01101" => level_vec_out <= "1011110001111111001100011111101111100011111011111101001110011111110111001110111001111011111111110101";
                    when "01110" => level_vec_out <= "1011110001111111001100011111101111100011111011111101001110011111110111001110111001111011111111110101";
                    when "01111" => level_vec_out <= "1011110001111111001101011111101111110011111111111101011110011111110111011110111001111011111111110101";
                    when "10000" => level_vec_out <= "1111110011111111001101011111101111110011111111111101011110011111110111011110111101111011111111110101";
                    when "10001" => level_vec_out <= "1111110111111111001101111111101111110011111111111101011110011111110111011110111101111011111111110101";
                    when "10010" => level_vec_out <= "1111110111111111001101111111101111110011111111111101011110011111110111011110111101111011111111110101";
                    when "10011" => level_vec_out <= "1111110111111111001101111111101111110011111111111101011110011111110111011110111101111011111111110101";
                    when "10100" => level_vec_out <= "1111110111111111001101111111111111110011111111111101011110111111110111011110111101111011111111110101";
                    when "10101" => level_vec_out <= "1111110111111111001101111111111111110011111111111101111111111111111111011111111101111011111111110101";
                    when "10110" => level_vec_out <= "1111110111111111001101111111111111111011111111111101111111111111111111011111111101111011111111110101";
                    when "10111" => level_vec_out <= "1111110111111111001101111111111111111011111111111111111111111111111111011111111111111111111111110101";
                    when "11000" => level_vec_out <= "1111110111111111001101111111111111111011111111111111111111111111111111011111111111111111111111110101";
                    when "11001" => level_vec_out <= "1111110111111111001101111111111111111011111111111111111111111111111111011111111111111111111111110101";
                    when "11010" => level_vec_out <= "1111110111111111101101111111111111111111111111111111111111111111111111011111111111111111111111110101";
                    when "11011" => level_vec_out <= "1111111111111111101101111111111111111111111111111111111111111111111111011111111111111111111111110101";
                    when "11100" => level_vec_out <= "1111111111111111101101111111111111111111111111111111111111111111111111011111111111111111111111110101";
                    when "11101" => level_vec_out <= "1111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111110101";
                when others => null;
                end case;
            when "1001" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1001101110101110010110101110101101010101010011011111011000110100011001010100010000110010001101101010";
                    when "00001" => level_vec_out <= "1001101110101110010110101110101101010101010011011111111000110110011001010100010000110010001101101010";
                    when "00010" => level_vec_out <= "1001101110101110010110101110101101010101010011011111111000110110011001010100011000110011001101101010";
                    when "00011" => level_vec_out <= "1101111110101110010110101110101101010101010011011111111000110111011001110100011000110011001101101010";
                    when "00100" => level_vec_out <= "1101111110101110010111101110101101010101010011011111111000110111011001110100011010110011001101101010";
                    when "00101" => level_vec_out <= "1101111110101110110111101110101101010101010011011111111000110111011001110100011010110011001101111010";
                    when "00110" => level_vec_out <= "1101111110101110110111101110101101010101010011011111111100110111011001110100011010110011001101111010";
                    when "00111" => level_vec_out <= "1101111110101110110111101110101101010101010011011111111110110111011001110100011010110011001101111010";
                    when "01000" => level_vec_out <= "1101111110101110110111101110101101010101010011011111111110110111011001110100011110110011001101111010";
                    when "01001" => level_vec_out <= "1101111110101110110111101110101101010101010011011111111110110111011011110100011110110011001101111010";
                    when "01010" => level_vec_out <= "1101111110101110110111101110101101010101010011011111111110110111011011110100011110110011001101111010";
                    when "01011" => level_vec_out <= "1101111110101110110111101110101101010101010011011111111110110111011011110100011110110011001101111110";
                    when "01100" => level_vec_out <= "1101111110101110110111101110101101010101010111011111111110110111011111110100011110110011001101111110";
                    when "01101" => level_vec_out <= "1101111110101110110111111110101101010101010111111111111110110111011111110110011110110011001101111110";
                    when "01110" => level_vec_out <= "1101111110101110110111111110101101010101010111111111111110110111011111110110011111110011011101111110";
                    when "01111" => level_vec_out <= "1101111110101110110111111110111101010101010111111111111110110111011111110110011111110011011101111110";
                    when "10000" => level_vec_out <= "1101111110101110110111111110111101010101010111111111111110110111011111110110011111110011011101111110";
                    when "10001" => level_vec_out <= "1101111110101110110111111110111111011101010111111111111110110111011111110110011111110011011101111110";
                    when "10010" => level_vec_out <= "1101111111101110110111111110111111011101010111111111111110110111011111110110011111110111111101111110";
                    when "10011" => level_vec_out <= "1101111111101110110111111110111111011101010111111111111110110111111111110110011111111111111101111110";
                    when "10100" => level_vec_out <= "1101111111101110110111111110111111011101010111111111111110110111111111110110011111111111111101111110";
                    when "10101" => level_vec_out <= "1111111111101110110111111110111111011101010111111111111110110111111111110111011111111111111101111110";
                    when "10110" => level_vec_out <= "1111111111101110110111111110111111111101010111111111111110110111111111110111011111111111111101111110";
                    when "10111" => level_vec_out <= "1111111111101110110111111110111111111101010111111111111110110111111111110111011111111111111101111110";
                    when "11000" => level_vec_out <= "1111111111101110110111111110111111111101010111111111111110110111111111110111011111111111111111111111";
                    when "11001" => level_vec_out <= "1111111111111110110111111110111111111101010111111111111110110111111111110111011111111111111111111111";
                    when "11010" => level_vec_out <= "1111111111111110110111111110111111111111010111111111111110110111111111110111011111111111111111111111";
                    when "11011" => level_vec_out <= "1111111111111110110111111111111111111111110111111111111111110111111111110111011111111111111111111111";
                    when "11100" => level_vec_out <= "1111111111111110110111111111111111111111110111111111111111110111111111110111011111111111111111111111";
                    when "11101" => level_vec_out <= "1111111111111110110111111111111111111111110111111111111111110111111111110111011111111111111111111111";
                when others => null;
                end case;
            when others => null;
        end case;
    end process;
end Behavioral;