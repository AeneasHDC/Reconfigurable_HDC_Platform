/**
 * @file level_hvec_gen_hdl.hpp
 * @brief This script generates HDL code for generating high-dimensional LEVEL vectors.
 * It is a novel method; for more information, please refer to our paper.
 *
 * @author Saeid Jamili and Marco Angioli
 * @note Author names are listed in alphabetical order.
 * @email <saeid.jamili@uniroma1.it>
 * @email <marco.angioli@uniroma1.it>
 *
 * @contributors
 *
 * @date Created: 24th July 2023
 * @date Last Updated: 23th August 2023
 *
 * @version 1.0.0
 *
 * @institute Sapienza University of Rome
 * @cite https://doi.org/10.xxxx/yyyyy
 *
 * @section DEPENDENCIES
 * - Dependency1: Description or version details.
 * - Dependency2: Description or version details.
 *
 * @section LICENSE
 * This file is part of the Aeneas HyperCompute Platform.
 *
 * Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 *
 * @section CHANGELOG
 * @version 1.0.0-dev - 23th August 2023
 * - Initial release
 *
 * @todo
 * - Complete level vector generator function
 * - Add training
 *
 * @see
 * -
 * -
 * -
 *
 */

module level_vec_gen (
    output reg [63:0] level_vec_out,
    input [2:0] frame_index,
    input [4:0] frame_id
);
    always @(*) begin
        // Update this function to match your requirements
        case (frame_index)
            0: begin
                case (frame_id)
                    0: level_vec_out = 64'b1110100110111100001011010111110100011111010000010010010001111111;
                    1: level_vec_out = 64'b1110100110111110011011110111110100011111010000010010010001111111;
                    2: level_vec_out = 64'b1110100110111110011011110111110100011111010000010110010001111111;
                    3: level_vec_out = 64'b1110100110111110011111110111110100011111010000010111010001111111;
                    4: level_vec_out = 64'b1110100110111110011111110111110100011111010000010111010001111111;
                    5: level_vec_out = 64'b1110100110111111011111110111111100011111010000010111010001111111;
                    6: level_vec_out = 64'b1110100110111111011111110111111100011111010000010111010011111111;
                    7: level_vec_out = 64'b1110100110111111011111110111111100111111010000010111010011111111;
                    8: level_vec_out = 64'b1110100110111111011111110111111100111111010000010111010011111111;
                    9: level_vec_out = 64'b1110100110111111011111110111111100111111010000010111010011111111;
                    10: level_vec_out = 64'b1110100110111111011111110111111100111111010000010111010011111111;
                    11: level_vec_out = 64'b1110100110111111011111110111111100111111010000010111010011111111;
                    12: level_vec_out = 64'b1110100110111111111111110111111100111111010000010111010011111111;
                    13: level_vec_out = 64'b1110100110111111111111110111111100111111010000010111010011111111;
                    14: level_vec_out = 64'b1110100110111111111111110111111100111111010000010111010111111111;
                    15: level_vec_out = 64'b1110100110111111111111110111111100111111010000010111010111111111;
                    16: level_vec_out = 64'b1110100110111111111111110111111101111111010000010111010111111111;
                    17: level_vec_out = 64'b1110100110111111111111110111111101111111010000010111010111111111;
                    18: level_vec_out = 64'b1110100110111111111111110111111101111111010000010111010111111111;
                    19: level_vec_out = 64'b1110100110111111111111110111111101111111110010010111010111111111;
                    20: level_vec_out = 64'b1110100110111111111111110111111101111111110010010111010111111111;
                    21: level_vec_out = 64'b1110100110111111111111110111111101111111110110010111010111111111;
                    22: level_vec_out = 64'b1110100110111111111111110111111101111111110110010111010111111111;
                    23: level_vec_out = 64'b1110100110111111111111110111111101111111110110010111010111111111;
                    24: level_vec_out = 64'b1110100110111111111111110111111101111111110110010111110111111111;
                    25: level_vec_out = 64'b1110101111111111111111110111111101111111110111010111110111111111;
                    26: level_vec_out = 64'b1110101111111111111111110111111101111111110111010111110111111111;
                    27: level_vec_out = 64'b1110101111111111111111110111111101111111110111010111110111111111;
                    28: level_vec_out = 64'b1110101111111111111111110111111111111111110111010111110111111111;
                    29: level_vec_out = 64'b1110101111111111111111111111111111111111110111010111110111111111;
                    30: level_vec_out = 64'b1111101111111111111111111111111111111111111111011111110111111111;
                    31: level_vec_out = 64'b1111101111111111111111111111111111111111111111111111110111111111;
                endcase
            end
            1: begin
                case (frame_id)
                    0: level_vec_out = 64'b1001000000101100111000110100010000111010010000001001111001100101;
                    1: level_vec_out = 64'b1001000000101100111000110100010000111010010000001001111001100101;
                    2: level_vec_out = 64'b1001000000101100111000110100010000111010010000001001111001100101;
                    3: level_vec_out = 64'b1001100000101100111000110100010000111010010001001001111001100101;
                    4: level_vec_out = 64'b1001100000101100111000110100011011111010010001001001111001101101;
                    5: level_vec_out = 64'b1001100000101101111000110100011011111010010001001001111001101101;
                    6: level_vec_out = 64'b1001100000101101111010110100011011111010010001001001111001101101;
                    7: level_vec_out = 64'b1001101000101101111010110100011011111010010001001001111011101101;
                    8: level_vec_out = 64'b1001101000101101111010110101011011111010010001001001111011101101;
                    9: level_vec_out = 64'b1001101011101101111010110101011011111010010001001001111011101101;
                    10: level_vec_out = 64'b1001101011101101111010110101011011111010010001001001111011101101;
                    11: level_vec_out = 64'b1001101011111101111010110101011011111010010001001001111011101101;
                    12: level_vec_out = 64'b1001101011111101111010111101011111111010010001001001111011101101;
                    13: level_vec_out = 64'b1001101011111101111010111101011111111010011001001001111011101101;
                    14: level_vec_out = 64'b1001101011111101111010111101011111111010011001001001111011101101;
                    15: level_vec_out = 64'b1001101011111101111010111101011111111010011001001101111011101101;
                    16: level_vec_out = 64'b1001101011111101111010111101011111111010011001001101111111101101;
                    17: level_vec_out = 64'b1001101011111101111010111101011111111110011001001101111111101101;
                    18: level_vec_out = 64'b1001101011111101111010111101011111111110011001001101111111101101;
                    19: level_vec_out = 64'b1001101011111101111010111101011111111110011001101111111111101101;
                    20: level_vec_out = 64'b1001111011111101111110111101011111111110011001101111111111101101;
                    21: level_vec_out = 64'b1001111011111101111110111101011111111110011001101111111111101101;
                    22: level_vec_out = 64'b1001111011111101111110111101011111111111011001101111111111101101;
                    23: level_vec_out = 64'b1001111011111101111110111101011111111111011001101111111111111101;
                    24: level_vec_out = 64'b1001111011111111111110111101011111111111111001101111111111111101;
                    25: level_vec_out = 64'b1001111111111111111111111101011111111111111001101111111111111101;
                    26: level_vec_out = 64'b1011111111111111111111111101011111111111111001101111111111111101;
                    27: level_vec_out = 64'b1011111111111111111111111101011111111111111001111111111111111101;
                    28: level_vec_out = 64'b1011111111111111111111111101011111111111111101111111111111111111;
                    29: level_vec_out = 64'b1111111111111111111111111101011111111111111101111111111111111111;
                    30: level_vec_out = 64'b1111111111111111111111111101011111111111111101111111111111111111;
                    31: level_vec_out = 64'b1111111111111111111111111101011111111111111101111111111111111111;
                endcase
            end
            2: begin
                case (frame_id)
                    0: level_vec_out = 64'b0001101010110101110101011110010011011100100110111000110101000011;
                    1: level_vec_out = 64'b0001101010110101110101011110010011011100100110111000110101000011;
                    2: level_vec_out = 64'b0001101010110101110101011110010011011100100110111000110101000011;
                    3: level_vec_out = 64'b1001101010110101110111011110010011011100100110111000110101000011;
                    4: level_vec_out = 64'b1001101010110101110111011110010011011100100110111000110101000011;
                    5: level_vec_out = 64'b1001101010110111111111011110010011011100100110111000110101000011;
                    6: level_vec_out = 64'b1001101010110111111111011110010011011100100110111100110101000011;
                    7: level_vec_out = 64'b1001101010110111111111011110010011011100100110111100110101010011;
                    8: level_vec_out = 64'b1001101010110111111111011110010011011100100110111101110101010011;
                    9: level_vec_out = 64'b1001111010110111111111011110010011011100100110111101110101010011;
                    10: level_vec_out = 64'b1001111010110111111111011110011011011100100110111101110101010011;
                    11: level_vec_out = 64'b1011111010111111111111011110011011011100100110111101110101010011;
                    12: level_vec_out = 64'b1011111010111111111111011110011011011100100110111101110101010011;
                    13: level_vec_out = 64'b1011111010111111111111011110011011011100100110111101111101010011;
                    14: level_vec_out = 64'b1011111010111111111111011110011011011100100110111101111101010011;
                    15: level_vec_out = 64'b1011111010111111111111011110011011011100100110111101111101010011;
                    16: level_vec_out = 64'b1011111110111111111111011110011011011100100111111101111101010011;
                    17: level_vec_out = 64'b1011111110111111111111011110011011011100100111111101111101110011;
                    18: level_vec_out = 64'b1011111110111111111111011110011011011100100111111101111101110011;
                    19: level_vec_out = 64'b1011111110111111111111011110011011011100100111111101111101110011;
                    20: level_vec_out = 64'b1011111110111111111111011110011011011100100111111101111101110011;
                    21: level_vec_out = 64'b1011111110111111111111011110011011011110100111111101111101110011;
                    22: level_vec_out = 64'b1011111110111111111111011110011011011110100111111101111101111011;
                    23: level_vec_out = 64'b1011111110111111111111011110011011011110100111111111111101111011;
                    24: level_vec_out = 64'b1011111110111111111111111110011011011110110111111111111101111011;
                    25: level_vec_out = 64'b1011111110111111111111111110111011011110110111111111111101111011;
                    26: level_vec_out = 64'b1011111110111111111111111110111011011110110111111111111111111011;
                    27: level_vec_out = 64'b1011111110111111111111111110111011111110111111111111111111111011;
                    28: level_vec_out = 64'b1011111110111111111111111110111111111110111111111111111111111011;
                    29: level_vec_out = 64'b1011111110111111111111111110111111111110111111111111111111111011;
                    30: level_vec_out = 64'b1111111110111111111111111111111111111110111111111111111111111011;
                    31: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                endcase
            end
            3: begin
                case (frame_id)
                    0: level_vec_out = 64'b1101101010001000101111010000001010110011110000110100001101110000;
                    1: level_vec_out = 64'b1101101010001000101111011000001010110011110000110100001101110000;
                    2: level_vec_out = 64'b1101101010001000101111011000001010110011110000110110001101110000;
                    3: level_vec_out = 64'b1101101010001000101111011000001010110011110001110110001101110000;
                    4: level_vec_out = 64'b1101101011001000101111011001001010110011110001110110001101110000;
                    5: level_vec_out = 64'b1101101011001000101111011001001010110011110001110110001111110000;
                    6: level_vec_out = 64'b1101101011001000101111011001001011110011110001110110001111110000;
                    7: level_vec_out = 64'b1101101011001000101111011001001111111011110001110110001111110000;
                    8: level_vec_out = 64'b1101101011011000101111011101001111111011110011110110001111110000;
                    9: level_vec_out = 64'b1101101011011000101111011101011111111011110011110110001111110000;
                    10: level_vec_out = 64'b1101101111011000111111011101011111111011110011110110001111110000;
                    11: level_vec_out = 64'b1101101111011000111111011101011111111011110011110110001111110000;
                    12: level_vec_out = 64'b1101101111011000111111011101011111111011110011110110001111110000;
                    13: level_vec_out = 64'b1101101111011000111111111101011111111011110011110110001111110010;
                    14: level_vec_out = 64'b1101101111011001111111111101011111111111110011110110001111110010;
                    15: level_vec_out = 64'b1101101111011101111111111101011111111111110011110110001111110010;
                    16: level_vec_out = 64'b1101111111011101111111111101011111111111110011110110001111111010;
                    17: level_vec_out = 64'b1111111111011101111111111101011111111111110011110110001111111010;
                    18: level_vec_out = 64'b1111111111111111111111111101111111111111110011110110001111111010;
                    19: level_vec_out = 64'b1111111111111111111111111111111111111111110011110110001111111010;
                    20: level_vec_out = 64'b1111111111111111111111111111111111111111110011110110001111111010;
                    21: level_vec_out = 64'b1111111111111111111111111111111111111111111011110110011111111010;
                    22: level_vec_out = 64'b1111111111111111111111111111111111111111111011110110011111111111;
                    23: level_vec_out = 64'b1111111111111111111111111111111111111111111011110110011111111111;
                    24: level_vec_out = 64'b1111111111111111111111111111111111111111111111110110011111111111;
                    25: level_vec_out = 64'b1111111111111111111111111111111111111111111111111110011111111111;
                    26: level_vec_out = 64'b1111111111111111111111111111111111111111111111111110011111111111;
                    27: level_vec_out = 64'b1111111111111111111111111111111111111111111111111110011111111111;
                    28: level_vec_out = 64'b1111111111111111111111111111111111111111111111111110011111111111;
                    29: level_vec_out = 64'b1111111111111111111111111111111111111111111111111110111111111111;
                    30: level_vec_out = 64'b1111111111111111111111111111111111111111111111111110111111111111;
                    31: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                endcase
            end
            4: begin
                case (frame_id)
                    0: level_vec_out = 64'b1110011111110101111100011001110100100011111110000110001101001111;
                    1: level_vec_out = 64'b1110011111110101111100011001110100100011111110001110001101001111;
                    2: level_vec_out = 64'b1110011111110101111100011001111100100011111110101110001101001111;
                    3: level_vec_out = 64'b1110011111110101111100011001111100100011111110101110001101001111;
                    4: level_vec_out = 64'b1110011111110101111100011001111100100011111110101110001101001111;
                    5: level_vec_out = 64'b1110011111110101111100011001111100100011111110101110011101001111;
                    6: level_vec_out = 64'b1110011111111101111100011001111100100011111110101110011101001111;
                    7: level_vec_out = 64'b1110011111111101111100011001111110100011111110101110011101001111;
                    8: level_vec_out = 64'b1110111111111101111100011001111110100011111110101110011101001111;
                    9: level_vec_out = 64'b1110111111111101111101011001111110110011111110101110011101001111;
                    10: level_vec_out = 64'b1110111111111101111101011001111110110011111110101111011101001111;
                    11: level_vec_out = 64'b1110111111111101111101011001111110110011111110101111011111001111;
                    12: level_vec_out = 64'b1110111111111101111101011101111110110011111110101111011111001111;
                    13: level_vec_out = 64'b1110111111111101111101011101111110110011111110101111011111001111;
                    14: level_vec_out = 64'b1110111111111101111101011101111110110011111110101111011111001111;
                    15: level_vec_out = 64'b1110111111111101111101011101111110110011111110101111011111001111;
                    16: level_vec_out = 64'b1110111111111101111101011101111110110011111110101111011111001111;
                    17: level_vec_out = 64'b1110111111111111111101011101111110110011111110101111011111001111;
                    18: level_vec_out = 64'b1110111111111111111101011101111110110011111110101111011111001111;
                    19: level_vec_out = 64'b1110111111111111111101011101111110110011111110101111011111001111;
                    20: level_vec_out = 64'b1110111111111111111101011101111110111011111110101111011111001111;
                    21: level_vec_out = 64'b1110111111111111111101011101111110111011111110101111011111001111;
                    22: level_vec_out = 64'b1110111111111111111101011101111110111011111111101111011111001111;
                    23: level_vec_out = 64'b1110111111111111111101011101111110111011111111101111011111101111;
                    24: level_vec_out = 64'b1110111111111111111101011101111110111011111111101111011111101111;
                    25: level_vec_out = 64'b1110111111111111111101011101111110111011111111101111011111101111;
                    26: level_vec_out = 64'b1110111111111111111101011111111110111011111111101111011111101111;
                    27: level_vec_out = 64'b1111111111111111111101011111111110111011111111101111011111101111;
                    28: level_vec_out = 64'b1111111111111111111111011111111110111011111111111111011111101111;
                    29: level_vec_out = 64'b1111111111111111111111011111111110111111111111111111011111101111;
                    30: level_vec_out = 64'b1111111111111111111111111111111110111111111111111111011111111111;
                    31: level_vec_out = 64'b1111111111111111111111111111111110111111111111111111111111111111;
                endcase
            end
            5: begin
                case (frame_id)
                    0: level_vec_out = 64'b1000001011010000011110011001101101000111100001100001000111101101;
                    1: level_vec_out = 64'b1000001011010000011110011001101101000111100001100001000111101101;
                    2: level_vec_out = 64'b1000101011010000011110011001101101000111100001100001000111101101;
                    3: level_vec_out = 64'b1000101011010000011110011001101101000111100001100001000111101101;
                    4: level_vec_out = 64'b1000101011010000011110011001101101000111100001100001000111101101;
                    5: level_vec_out = 64'b1000101011010000011110011001101101000111100001100001000111101101;
                    6: level_vec_out = 64'b1000101011010000011110011001101101000111100001100001000111101101;
                    7: level_vec_out = 64'b1000101011010000011110011001101101000111100001100001000111101101;
                    8: level_vec_out = 64'b1000101011010000011110011001101101000111110001100001000111101101;
                    9: level_vec_out = 64'b1000101011010000011110011001101101000111110001100001001111101101;
                    10: level_vec_out = 64'b1000101011010000011110011001101101000111110101100001001111101101;
                    11: level_vec_out = 64'b1000101011010000011110011001101101000111110101100001001111101101;
                    12: level_vec_out = 64'b1000101011010001011110011011101101000111110101100011001111101101;
                    13: level_vec_out = 64'b1000101011010001011110011011101101110111110101100011001111101101;
                    14: level_vec_out = 64'b1000101011110001111110011011101101110111110101100011001111101101;
                    15: level_vec_out = 64'b1100101011110001111110011011101101110111110101100111001111101101;
                    16: level_vec_out = 64'b1100101111110001111110011011101101110111110101100111001111101101;
                    17: level_vec_out = 64'b1100101111110001111110011011101101110111111101100111001111101111;
                    18: level_vec_out = 64'b1100101111110001111111011011101101110111111101100111011111101111;
                    19: level_vec_out = 64'b1100111111110001111111011011101101110111111101100111011111111111;
                    20: level_vec_out = 64'b1100111111110001111111011011101101110111111101110111011111111111;
                    21: level_vec_out = 64'b1100111111110001111111011011101101111111111101111111011111111111;
                    22: level_vec_out = 64'b1100111111110001111111011011101101111111111111111111011111111111;
                    23: level_vec_out = 64'b1100111111110101111111011011101101111111111111111111011111111111;
                    24: level_vec_out = 64'b1100111111110101111111011011101101111111111111111111011111111111;
                    25: level_vec_out = 64'b1100111111110101111111011011101101111111111111111111011111111111;
                    26: level_vec_out = 64'b1101111111111101111111011011101101111111111111111111011111111111;
                    27: level_vec_out = 64'b1101111111111111111111011111101101111111111111111111011111111111;
                    28: level_vec_out = 64'b1111111111111111111111011111101101111111111111111111111111111111;
                    29: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    30: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    31: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                endcase
            end
            6: begin
                case (frame_id)
                    0: level_vec_out = 64'b0011011001110000111110101010111100100010001111111000101100010001;
                    1: level_vec_out = 64'b0011011001110000111110101010111100100010001111111000111100010001;
                    2: level_vec_out = 64'b0011011001110000111110101010111100100010001111111000111110010001;
                    3: level_vec_out = 64'b0011011001110000111110101010111100100010001111111000111110010001;
                    4: level_vec_out = 64'b1011011001110000111110101010111100100010001111111000111110010001;
                    5: level_vec_out = 64'b1011011001110010111110101010111100100010001111111000111110010001;
                    6: level_vec_out = 64'b1111011001110110111110101010111100100010001111111000111110010001;
                    7: level_vec_out = 64'b1111011001110110111110101010111100100010001111111000111110010001;
                    8: level_vec_out = 64'b1111011001110110111110101010111100100010001111111000111110010001;
                    9: level_vec_out = 64'b1111011001110110111110101010111100100010001111111000111110010001;
                    10: level_vec_out = 64'b1111011001110110111110101010111100100010001111111000111110010001;
                    11: level_vec_out = 64'b1111011011110110111110101010111100100010001111111000111110010101;
                    12: level_vec_out = 64'b1111011011110111111110101010111100100010001111111000111110010101;
                    13: level_vec_out = 64'b1111011011110111111110101010111100100010001111111000111110010101;
                    14: level_vec_out = 64'b1111011011110111111110101010111100100010001111111010111110011101;
                    15: level_vec_out = 64'b1111011011110111111110101010111110100010001111111010111110011101;
                    16: level_vec_out = 64'b1111011011110111111110101010111110100010001111111010111110111101;
                    17: level_vec_out = 64'b1111011111110111111110101010111110100010001111111110111110111101;
                    18: level_vec_out = 64'b1111011111110111111110101010111110100010001111111110111110111101;
                    19: level_vec_out = 64'b1111011111110111111110101010111110110010001111111110111110111101;
                    20: level_vec_out = 64'b1111011111111111111110101010111111110010001111111110111110111111;
                    21: level_vec_out = 64'b1111011111111111111110101010111111110010011111111110111110111111;
                    22: level_vec_out = 64'b1111011111111111111110101010111111110010011111111111111110111111;
                    23: level_vec_out = 64'b1111011111111111111110101010111111110010011111111111111110111111;
                    24: level_vec_out = 64'b1111011111111111111110101010111111110010111111111111111110111111;
                    25: level_vec_out = 64'b1111111111111111111110101010111111110010111111111111111110111111;
                    26: level_vec_out = 64'b1111111111111111111110111011111111110010111111111111111110111111;
                    27: level_vec_out = 64'b1111111111111111111110111011111111110110111111111111111111111111;
                    28: level_vec_out = 64'b1111111111111111111110111011111111110110111111111111111111111111;
                    29: level_vec_out = 64'b1111111111111111111110111011111111110110111111111111111111111111;
                    30: level_vec_out = 64'b1111111111111111111110111011111111110111111111111111111111111111;
                    31: level_vec_out = 64'b1111111111111111111111111011111111111111111111111111111111111111;
                endcase
            end
            7: begin
                case (frame_id)
                    0: level_vec_out = 64'b1010101000111001011010110100000011011100001100111000001001100011;
                    1: level_vec_out = 64'b1010101000111001011010110100000011011100001111111000001001100011;
                    2: level_vec_out = 64'b1010101000111001111010110100000011011100001111111010001001100011;
                    3: level_vec_out = 64'b1010101000111001111010110110000011011100001111111010001001100011;
                    4: level_vec_out = 64'b1010101000111001111010110110000111011100001111111010001001100011;
                    5: level_vec_out = 64'b1010101000111001111010110110000111011100001111111010001001100011;
                    6: level_vec_out = 64'b1010101000111001111010110110000111011110001111111010001001100011;
                    7: level_vec_out = 64'b1010101000111101111010110110000111011110001111111010001001100011;
                    8: level_vec_out = 64'b1010111000111101111010110110000111011110001111111010001001100011;
                    9: level_vec_out = 64'b1010111000111101111010110110000111011110011111111010001001100011;
                    10: level_vec_out = 64'b1010111100111101111010110110100111011110011111111110001001100011;
                    11: level_vec_out = 64'b1010111100111101111110110110100111011110011111111110001001100111;
                    12: level_vec_out = 64'b1010111100111101111110110110100111011110011111111110001001100111;
                    13: level_vec_out = 64'b1010111100111101111110110110101111011110011111111110101001100111;
                    14: level_vec_out = 64'b1110111100111101111110110110101111011110011111111110101001100111;
                    15: level_vec_out = 64'b1110111100111101111110110110111111011111011111111110111001100111;
                    16: level_vec_out = 64'b1110111100111101111110110110111111011111011111111110111001100111;
                    17: level_vec_out = 64'b1110111100111101111110110110111111011111011111111110111001100111;
                    18: level_vec_out = 64'b1110111100111111111110110110111111011111011111111110111001111111;
                    19: level_vec_out = 64'b1110111100111111111110110110111111011111011111111110111001111111;
                    20: level_vec_out = 64'b1110111100111111111110110110111111011111011111111110111011111111;
                    21: level_vec_out = 64'b1110111101111111111110110110111111011111011111111110111011111111;
                    22: level_vec_out = 64'b1110111101111111111110110110111111011111111111111110111011111111;
                    23: level_vec_out = 64'b1111111111111111111110111111111111011111111111111110111011111111;
                    24: level_vec_out = 64'b1111111111111111111110111111111111011111111111111111111011111111;
                    25: level_vec_out = 64'b1111111111111111111110111111111111011111111111111111111011111111;
                    26: level_vec_out = 64'b1111111111111111111110111111111111111111111111111111111011111111;
                    27: level_vec_out = 64'b1111111111111111111110111111111111111111111111111111111011111111;
                    28: level_vec_out = 64'b1111111111111111111110111111111111111111111111111111111011111111;
                    29: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111011111111;
                    30: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111011111111;
                    31: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111011111111;
                endcase
            end
        endcase
    end
endmodule