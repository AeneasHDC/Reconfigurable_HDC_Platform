/**
 * @file level_hvec_gen_hdl.hpp
 * @brief This script generates HDL code for generating high-dimensional LEVEL vectors.
 * It is a novel method; for more information, please refer to our paper.
 *
 * @author Saeid Jamili and Marco Angioli
 * @note Author names are listed in alphabetical order.
 * @email <saeid.jamili@uniroma1.it>
 * @email <marco.angioli@uniroma1.it>
 *
 * @contributors
 *
 * @date Created: 24th July 2023
 * @date Last Updated: 23th August 2023
 *
 * @version 1.0.0
 *
 * @institute Sapienza University of Rome
 * @cite https://doi.org/10.xxxx/yyyyy
 *
 * @section DEPENDENCIES
 * - Dependency1: Description or version details.
 * - Dependency2: Description or version details.
 *
 * @section LICENSE
 * This file is part of the Aeneas HyperCompute Platform.
 *
 * Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 *
 * @section CHANGELOG
 * @version 1.0.0-dev - 23th August 2023
 * - Initial release
 *
 * @todo
 * - Complete level vector generator function
 * - Add training
 *
 * @see
 * -
 * -
 * -
 *
 */

module level_vec_gen (
    output reg [63:0] level_vec_out,
    input [2:0] frame_index,
    input [4:0] frame_id
);
    always @(*) begin
        // Update this function to match your requirements
        case (frame_index)
            0: begin
                case (frame_id)
                    0: level_vec_out = 64'b1111100011110101011011110101100111100000010100101000101000110000;
                    1: level_vec_out = 64'b1111100011110101011011110101100111100000010100101000101000110000;
                    2: level_vec_out = 64'b1111101011110101011011110101100111100000010100101000101000110000;
                    3: level_vec_out = 64'b1111101011110101011011110101100111100000010100101000101000110000;
                    4: level_vec_out = 64'b1111101011110101011011110101100111100000010100101000101000110000;
                    5: level_vec_out = 64'b1111101011111101011011110101100111100010010100101000101000110000;
                    6: level_vec_out = 64'b1111101011111101011011110101100111100010010101101000101000110000;
                    7: level_vec_out = 64'b1111101011111101011011110101100111100010011101101000101000110000;
                    8: level_vec_out = 64'b1111101011111101011011110101100111100010011101101000101000110000;
                    9: level_vec_out = 64'b1111101011111101011011110101110111100010011101101000101000110000;
                    10: level_vec_out = 64'b1111101011111101011011110101111111100011111101101000101000110000;
                    11: level_vec_out = 64'b1111101011111101011011110101111111100011111101101000111000110001;
                    12: level_vec_out = 64'b1111101011111101011111110101111111100011111101101000111000110001;
                    13: level_vec_out = 64'b1111101011111101011111110101111111100011111101101000111000110001;
                    14: level_vec_out = 64'b1111101011111101011111110101111111100011111101101000111000111011;
                    15: level_vec_out = 64'b1111101011111101011111110101111111100011111101101000111100111011;
                    16: level_vec_out = 64'b1111101011111101011111110101111111100011111101101000111100111011;
                    17: level_vec_out = 64'b1111101011111111011111110101111111100011111101101000111100111011;
                    18: level_vec_out = 64'b1111101011111111011111110101111111100011111101101000111100111011;
                    19: level_vec_out = 64'b1111101011111111011111110101111111100011111101101001111100111011;
                    20: level_vec_out = 64'b1111101011111111011111110101111111100011111101101001111101111011;
                    21: level_vec_out = 64'b1111101011111111011111110101111111111011111101101101111101111011;
                    22: level_vec_out = 64'b1111101011111111011111110101111111111011111101101101111101111111;
                    23: level_vec_out = 64'b1111101011111111011111110101111111111011111101101101111101111111;
                    24: level_vec_out = 64'b1111101011111111011111111101111111111111111101101101111101111111;
                    25: level_vec_out = 64'b1111101011111111011111111101111111111111111101101101111101111111;
                    26: level_vec_out = 64'b1111101011111111011111111101111111111111111101111101111101111111;
                    27: level_vec_out = 64'b1111101011111111111111111101111111111111111101111101111101111111;
                    28: level_vec_out = 64'b1111101011111111111111111101111111111111111101111101111111111111;
                    29: level_vec_out = 64'b1111101011111111111111111111111111111111111101111101111111111111;
                    30: level_vec_out = 64'b1111111011111111111111111111111111111111111101111101111111111111;
                    31: level_vec_out = 64'b1111111011111111111111111111111111111111111101111111111111111111;
                endcase
            end
            1: begin
                case (frame_id)
                    0: level_vec_out = 64'b1010100001101100010010010010110000011001000010000000001111011111;
                    1: level_vec_out = 64'b1010100001101100010010010010110000011001000010100000001111011111;
                    2: level_vec_out = 64'b1010100001101100010011010010110000011001000010100000001111011111;
                    3: level_vec_out = 64'b1010100001101100010111010010110000011001000010100000001111011111;
                    4: level_vec_out = 64'b1110100001101110010111010010110000011001001010100000001111011111;
                    5: level_vec_out = 64'b1110100101101111010111010010110100011001001010100000001111011111;
                    6: level_vec_out = 64'b1110100101101111010111010010110100011001001010100000101111011111;
                    7: level_vec_out = 64'b1110100101101111010111010010110100011001001010100000101111011111;
                    8: level_vec_out = 64'b1110100101101111011111010010110100011001001010100000101111011111;
                    9: level_vec_out = 64'b1110100101101111011111010010111100011001001010100000101111011111;
                    10: level_vec_out = 64'b1110100101101111011111010010111100011001001010100010101111011111;
                    11: level_vec_out = 64'b1110100101101111011111010010111100011001001010100011101111011111;
                    12: level_vec_out = 64'b1110100111101111011111010011111100011001001010100011101111011111;
                    13: level_vec_out = 64'b1110100111101111011111010011111100011001011010110011101111011111;
                    14: level_vec_out = 64'b1110100111101111011111010011111100011001011010110011101111011111;
                    15: level_vec_out = 64'b1110100111101111011111010011111100011001011010110011101111011111;
                    16: level_vec_out = 64'b1110100111101111011111010011111100011011011010110111101111011111;
                    17: level_vec_out = 64'b1110100111101111011111010011111100011011011010110111101111011111;
                    18: level_vec_out = 64'b1110101111101111011111010011111100011011011011110111111111011111;
                    19: level_vec_out = 64'b1110101111101111011111010011111100011011011011110111111111011111;
                    20: level_vec_out = 64'b1110101111101111111111010111111100011011011011110111111111011111;
                    21: level_vec_out = 64'b1110101111111111111111010111111100011011011111111111111111011111;
                    22: level_vec_out = 64'b1110101111111111111111011111111100011011011111111111111111011111;
                    23: level_vec_out = 64'b1111101111111111111111011111111100011011011111111111111111011111;
                    24: level_vec_out = 64'b1111101111111111111111011111111100111011011111111111111111011111;
                    25: level_vec_out = 64'b1111101111111111111111011111111100111011011111111111111111111111;
                    26: level_vec_out = 64'b1111111111111111111111011111111100111011011111111111111111111111;
                    27: level_vec_out = 64'b1111111111111111111111011111111100111111011111111111111111111111;
                    28: level_vec_out = 64'b1111111111111111111111011111111101111111011111111111111111111111;
                    29: level_vec_out = 64'b1111111111111111111111111111111111111111011111111111111111111111;
                    30: level_vec_out = 64'b1111111111111111111111111111111111111111011111111111111111111111;
                    31: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                endcase
            end
            2: begin
                case (frame_id)
                    0: level_vec_out = 64'b0000010100010110010111010110110110001110110100010110110110010100;
                    1: level_vec_out = 64'b0000010100010110010111010110110110001110110110010110110110010100;
                    2: level_vec_out = 64'b0000010100010110010111010110110110001110110110010110110110010100;
                    3: level_vec_out = 64'b0000010100010110011111010110110110001110110110010110110110010100;
                    4: level_vec_out = 64'b0100010100010110011111010110110110001110110110010110110110010110;
                    5: level_vec_out = 64'b0100010100010110011111010110110110001110110110010110110110010110;
                    6: level_vec_out = 64'b0100010100010110011111010110110110001110110110011110110110010110;
                    7: level_vec_out = 64'b0100010100010111011111010110110110001110110110011110110110010110;
                    8: level_vec_out = 64'b0100010100010111011111011110110111001110110110011110110110010110;
                    9: level_vec_out = 64'b0100010100010111011111011110110111001110110111011110110110010110;
                    10: level_vec_out = 64'b0100010100010111011111011110110111001110110111011110110110010110;
                    11: level_vec_out = 64'b0100010100010111011111011110110111001110110111011110110110010111;
                    12: level_vec_out = 64'b0100010100010111011111011110110111001110110111011110110110010111;
                    13: level_vec_out = 64'b0100010100010111111111011110110111101110110111011110110110010111;
                    14: level_vec_out = 64'b0100010100010111111111011110110111101110110111011110110111010111;
                    15: level_vec_out = 64'b0110010100010111111111011110110111101111110111011110110111010111;
                    16: level_vec_out = 64'b0110010100010111111111111110110111101111110111011110110111010111;
                    17: level_vec_out = 64'b0110010100010111111111111110110111111111110111011110110111010111;
                    18: level_vec_out = 64'b0110010100010111111111111111110111111111110111011110110111010111;
                    19: level_vec_out = 64'b0110010100010111111111111111110111111111110111011110110111110111;
                    20: level_vec_out = 64'b0110010100010111111111111111110111111111110111011110110111110111;
                    21: level_vec_out = 64'b0110010100010111111111111111110111111111110111011110110111110111;
                    22: level_vec_out = 64'b0110010100010111111111111111110111111111110111011110110111110111;
                    23: level_vec_out = 64'b1110010100010111111111111111110111111111110111011110110111110111;
                    24: level_vec_out = 64'b1110010100010111111111111111110111111111110111111110110111110111;
                    25: level_vec_out = 64'b1110010100010111111111111111110111111111111111111111110111110111;
                    26: level_vec_out = 64'b1110010100010111111111111111110111111111111111111111110111110111;
                    27: level_vec_out = 64'b1110111100010111111111111111110111111111111111111111110111110111;
                    28: level_vec_out = 64'b1111111100011111111111111111110111111111111111111111110111110111;
                    29: level_vec_out = 64'b1111111100011111111111111111110111111111111111111111110111110111;
                    30: level_vec_out = 64'b1111111110111111111111111111110111111111111111111111110111110111;
                    31: level_vec_out = 64'b1111111110111111111111111111111111111111111111111111110111111111;
                endcase
            end
            3: begin
                case (frame_id)
                    0: level_vec_out = 64'b1011111001111111101000100111010001101100001001011000010000111110;
                    1: level_vec_out = 64'b1011111001111111111000100111010001101100101001011000010000111110;
                    2: level_vec_out = 64'b1011111001111111111000100111010001101100101001011000010000111110;
                    3: level_vec_out = 64'b1011111001111111111000100111010001101100101011011000010000111110;
                    4: level_vec_out = 64'b1011111001111111111000100111010001101100101011011000010000111110;
                    5: level_vec_out = 64'b1011111001111111111001100111010001101100101011011000010011111110;
                    6: level_vec_out = 64'b1011111001111111111001100111110001101100101011011000010011111110;
                    7: level_vec_out = 64'b1011111101111111111011100111110101101100101011011000010011111110;
                    8: level_vec_out = 64'b1011111101111111111011100111110101101110101011011101010011111110;
                    9: level_vec_out = 64'b1111111101111111111011100111110101101110101011011101010011111110;
                    10: level_vec_out = 64'b1111111111111111111011100111110101101110101011011101010111111110;
                    11: level_vec_out = 64'b1111111111111111111011100111110101101110101011011101010111111110;
                    12: level_vec_out = 64'b1111111111111111111011100111110101101110101011011101110111111110;
                    13: level_vec_out = 64'b1111111111111111111011100111110101101110101011011101110111111111;
                    14: level_vec_out = 64'b1111111111111111111011100111110101101110101111011101110111111111;
                    15: level_vec_out = 64'b1111111111111111111011100111110101101110101111011101110111111111;
                    16: level_vec_out = 64'b1111111111111111111011100111110101101110101111011101110111111111;
                    17: level_vec_out = 64'b1111111111111111111011100111110101101110101111011101110111111111;
                    18: level_vec_out = 64'b1111111111111111111011100111110101101110101111011101110111111111;
                    19: level_vec_out = 64'b1111111111111111111011100111110111101110101111011101110111111111;
                    20: level_vec_out = 64'b1111111111111111111011100111110111101110101111011101111111111111;
                    21: level_vec_out = 64'b1111111111111111111011100111110111101110101111011101111111111111;
                    22: level_vec_out = 64'b1111111111111111111011100111110111101110101111011101111111111111;
                    23: level_vec_out = 64'b1111111111111111111011110111110111101110101111011101111111111111;
                    24: level_vec_out = 64'b1111111111111111111011111111110111101110101111011101111111111111;
                    25: level_vec_out = 64'b1111111111111111111011111111110111101110111111011101111111111111;
                    26: level_vec_out = 64'b1111111111111111111011111111111111101111111111011111111111111111;
                    27: level_vec_out = 64'b1111111111111111111011111111111111101111111111011111111111111111;
                    28: level_vec_out = 64'b1111111111111111111011111111111111101111111111111111111111111111;
                    29: level_vec_out = 64'b1111111111111111111011111111111111101111111111111111111111111111;
                    30: level_vec_out = 64'b1111111111111111111011111111111111111111111111111111111111111111;
                    31: level_vec_out = 64'b1111111111111111111011111111111111111111111111111111111111111111;
                endcase
            end
            4: begin
                case (frame_id)
                    0: level_vec_out = 64'b1001110001111110111000000100000111101110110001010111010010010100;
                    1: level_vec_out = 64'b1001110001111110111000000110000111101110110001110111010010010100;
                    2: level_vec_out = 64'b1001110001111110111000000110000111101110110001110111010010010100;
                    3: level_vec_out = 64'b1011110001111110111000000110000111101110110001110111010010010100;
                    4: level_vec_out = 64'b1011110001111110111000000110000111101110110001110111010010010100;
                    5: level_vec_out = 64'b1011110001111110111000000110000111101110110001110111010010010100;
                    6: level_vec_out = 64'b1111110001111110111000000111000111101110110001110111010010010100;
                    7: level_vec_out = 64'b1111110001111110111000000111000111101110111001110111010010010100;
                    8: level_vec_out = 64'b1111110001111110111000000111000111101110111001110111010010010100;
                    9: level_vec_out = 64'b1111110001111110111000000111000111101110111001110111010010010100;
                    10: level_vec_out = 64'b1111110001111110111000000111000111101110111001110111010010010100;
                    11: level_vec_out = 64'b1111110001111110111000000111000111101110111001110111010010010100;
                    12: level_vec_out = 64'b1111110001111110111000000111000111101110111001110111010010010100;
                    13: level_vec_out = 64'b1111110001111110111000000111000111101110111001110111010010010100;
                    14: level_vec_out = 64'b1111110001111110111001000111000111101110111001111111010010010100;
                    15: level_vec_out = 64'b1111110001111110111001101111000111101110111001111111010011110100;
                    16: level_vec_out = 64'b1111110001111110111001101111010111101110111001111111010011110100;
                    17: level_vec_out = 64'b1111110001111110111001101111010111101110111011111111011011110100;
                    18: level_vec_out = 64'b1111110001111110111011101111010111101110111111111111011111110100;
                    19: level_vec_out = 64'b1111110001111111111011101111010111101111111111111111011111110100;
                    20: level_vec_out = 64'b1111110001111111111111101111011111101111111111111111011111110100;
                    21: level_vec_out = 64'b1111110001111111111111101111011111101111111111111111011111110100;
                    22: level_vec_out = 64'b1111111011111111111111111111011111101111111111111111011111110100;
                    23: level_vec_out = 64'b1111111011111111111111111111011111101111111111111111011111111100;
                    24: level_vec_out = 64'b1111111011111111111111111111111111101111111111111111011111111101;
                    25: level_vec_out = 64'b1111111011111111111111111111111111101111111111111111011111111101;
                    26: level_vec_out = 64'b1111111011111111111111111111111111101111111111111111011111111111;
                    27: level_vec_out = 64'b1111111011111111111111111111111111111111111111111111011111111111;
                    28: level_vec_out = 64'b1111111011111111111111111111111111111111111111111111111111111111;
                    29: level_vec_out = 64'b1111111011111111111111111111111111111111111111111111111111111111;
                    30: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    31: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                endcase
            end
            5: begin
                case (frame_id)
                    0: level_vec_out = 64'b0101011101100111110101010111110110100111100011111010101010101111;
                    1: level_vec_out = 64'b0101011101100111110101010111110110100111100011111010101010101111;
                    2: level_vec_out = 64'b0101011101100111110111010111110110100111100011111010101010101111;
                    3: level_vec_out = 64'b0101011101100111110111010111110110100111100011111011101011101111;
                    4: level_vec_out = 64'b1101011101100111110111010111110111100111100011111011101011101111;
                    5: level_vec_out = 64'b1101011101100111110111010111110111100111100011111011101011101111;
                    6: level_vec_out = 64'b1101011101100111110111010111110111100111100011111011101011101111;
                    7: level_vec_out = 64'b1101011101100111110111010111110111100111100011111011101011101111;
                    8: level_vec_out = 64'b1101011101100111110111010111110111100111100011111011101011101111;
                    9: level_vec_out = 64'b1101011101100111110111010111110111100111100011111011101011101111;
                    10: level_vec_out = 64'b1101011101100111110111010111110111100111110011111011101011101111;
                    11: level_vec_out = 64'b1101011101100111111111010111110111100111110011111011111011101111;
                    12: level_vec_out = 64'b1101011101100111111111110111110111101111110011111111111011101111;
                    13: level_vec_out = 64'b1101011101100111111111110111110111101111110011111111111011101111;
                    14: level_vec_out = 64'b1101011101100111111111110111110111101111110011111111111011101111;
                    15: level_vec_out = 64'b1101011101100111111111110111110111101111110011111111111011101111;
                    16: level_vec_out = 64'b1101111101101111111111110111110111101111110011111111111011101111;
                    17: level_vec_out = 64'b1101111101101111111111110111110111101111110011111111111011101111;
                    18: level_vec_out = 64'b1101111101101111111111110111110111101111110011111111111011101111;
                    19: level_vec_out = 64'b1101111101101111111111110111110111101111110111111111111011101111;
                    20: level_vec_out = 64'b1101111101101111111111110111110111101111110111111111111011101111;
                    21: level_vec_out = 64'b1101111101101111111111110111110111101111110111111111111011101111;
                    22: level_vec_out = 64'b1101111101101111111111110111110111101111110111111111111011111111;
                    23: level_vec_out = 64'b1101111101101111111111110111110111101111110111111111111011111111;
                    24: level_vec_out = 64'b1101111101101111111111111111110111101111110111111111111011111111;
                    25: level_vec_out = 64'b1101111101101111111111111111110111101111110111111111111011111111;
                    26: level_vec_out = 64'b1101111101111111111111111111110111101111110111111111111011111111;
                    27: level_vec_out = 64'b1101111101111111111111111111110111111111110111111111111011111111;
                    28: level_vec_out = 64'b1101111101111111111111111111110111111111110111111111111011111111;
                    29: level_vec_out = 64'b1101111111111111111111111111110111111111111111111111111011111111;
                    30: level_vec_out = 64'b1111111111111111111111111111110111111111111111111111111011111111;
                    31: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                endcase
            end
            6: begin
                case (frame_id)
                    0: level_vec_out = 64'b0110000011000110001100101111110000100110001101001010100100000001;
                    1: level_vec_out = 64'b0110000011000110001100101111110000100110101101001010100100000001;
                    2: level_vec_out = 64'b0111000011001110001100101111110000100110101101001010100100000001;
                    3: level_vec_out = 64'b0111000011001110001100101111110001100110101101001010100100000001;
                    4: level_vec_out = 64'b0111000011001110001100101111110001100110101101001010100100000001;
                    5: level_vec_out = 64'b0111000011001110001100101111110001100110101101001010100100000001;
                    6: level_vec_out = 64'b0111000111001110001100101111110001100110101101001010100100000001;
                    7: level_vec_out = 64'b0111000111001110001100101111110001100110101101001010110101000001;
                    8: level_vec_out = 64'b0111000111001110001100101111110001100110101101001010110101000001;
                    9: level_vec_out = 64'b0111000111001110001100101111110011100110101101001010110101000001;
                    10: level_vec_out = 64'b0111000111001110001100101111110011100110101101001110110101000001;
                    11: level_vec_out = 64'b0111011111001110001100101111110011100110101101001110110101000001;
                    12: level_vec_out = 64'b0111011111001110001100101111110111100110101101001110110101000001;
                    13: level_vec_out = 64'b1111011111001110001100101111111111100110101101001110110101000001;
                    14: level_vec_out = 64'b1111011111001110001100101111111111100110101101001110110101000011;
                    15: level_vec_out = 64'b1111011111001110001100101111111111100110101101001110110101000011;
                    16: level_vec_out = 64'b1111011111001110001101101111111111100110101101001110110101000011;
                    17: level_vec_out = 64'b1111011111001110001101101111111111100110101101001110111101000111;
                    18: level_vec_out = 64'b1111011111001110001101101111111111100110101101001110111101000111;
                    19: level_vec_out = 64'b1111011111011110001101101111111111100110101101001110111101000111;
                    20: level_vec_out = 64'b1111011111111110001101101111111111100110111101001110111101000111;
                    21: level_vec_out = 64'b1111011111111110001101101111111111101110111101001110111101000111;
                    22: level_vec_out = 64'b1111011111111110001101101111111111101110111101001110111101001111;
                    23: level_vec_out = 64'b1111011111111110111101101111111111101110111101001111111101001111;
                    24: level_vec_out = 64'b1111011111111110111101101111111111101110111101001111111101001111;
                    25: level_vec_out = 64'b1111011111111111111101101111111111111110111111001111111101001111;
                    26: level_vec_out = 64'b1111111111111111111101101111111111111110111111001111111101001111;
                    27: level_vec_out = 64'b1111111111111111111101111111111111111110111111011111111101001111;
                    28: level_vec_out = 64'b1111111111111111111101111111111111111110111111011111111101101111;
                    29: level_vec_out = 64'b1111111111111111111101111111111111111110111111111111111101111111;
                    30: level_vec_out = 64'b1111111111111111111111111111111111111110111111111111111101111111;
                    31: level_vec_out = 64'b1111111111111111111111111111111111111110111111111111111101111111;
                endcase
            end
            7: begin
                case (frame_id)
                    0: level_vec_out = 64'b1110010101010110011111010001010100111000101001111110100011001010;
                    1: level_vec_out = 64'b1110010101010110011111010001010100111000101001111110110011001010;
                    2: level_vec_out = 64'b1110010101010110011111010011010100111010111001111110110011001010;
                    3: level_vec_out = 64'b1110010101010110011111010011010100111010111011111110110011001010;
                    4: level_vec_out = 64'b1110010101010110011111010011010100111110111011111110110011001010;
                    5: level_vec_out = 64'b1110010101010110011111010011010100111110111011111110110011001010;
                    6: level_vec_out = 64'b1110010101010110011111010011010100111110111011111110111011001010;
                    7: level_vec_out = 64'b1110010101010110011111010011010100111110111011111110111011001010;
                    8: level_vec_out = 64'b1110011101011110011111010011010100111110111011111110111011001010;
                    9: level_vec_out = 64'b1110011101011111011111010111010100111111111011111110111011001010;
                    10: level_vec_out = 64'b1110011101011111011111010111010100111111111011111110111011001010;
                    11: level_vec_out = 64'b1110011101011111011111010111010100111111111011111110111011001010;
                    12: level_vec_out = 64'b1110011101011111011111010111010100111111111011111110111011001010;
                    13: level_vec_out = 64'b1110011101011111011111010111010100111111111011111110111011011010;
                    14: level_vec_out = 64'b1110011101011111011111010111010100111111111011111110111111011010;
                    15: level_vec_out = 64'b1110011101011111011111010111010100111111111011111110111111111010;
                    16: level_vec_out = 64'b1110111101011111011111010111010100111111111011111110111111111010;
                    17: level_vec_out = 64'b1110111101011111011111010111011110111111111011111110111111111010;
                    18: level_vec_out = 64'b1110111101011111111111010111011110111111111011111110111111111010;
                    19: level_vec_out = 64'b1110111101011111111111010111011110111111111011111111111111111010;
                    20: level_vec_out = 64'b1110111101011111111111010111011110111111111011111111111111111010;
                    21: level_vec_out = 64'b1111111101011111111111010111011110111111111011111111111111111010;
                    22: level_vec_out = 64'b1111111101011111111111010111111110111111111011111111111111111010;
                    23: level_vec_out = 64'b1111111101011111111111010111111111111111111011111111111111111010;
                    24: level_vec_out = 64'b1111111101011111111111010111111111111111111011111111111111111010;
                    25: level_vec_out = 64'b1111111101011111111111010111111111111111111011111111111111111011;
                    26: level_vec_out = 64'b1111111101011111111111010111111111111111111011111111111111111011;
                    27: level_vec_out = 64'b1111111101011111111111010111111111111111111011111111111111111011;
                    28: level_vec_out = 64'b1111111101011111111111010111111111111111111111111111111111111011;
                    29: level_vec_out = 64'b1111111101011111111111110111111111111111111111111111111111111011;
                    30: level_vec_out = 64'b1111111111011111111111110111111111111111111111111111111111111011;
                    31: level_vec_out = 64'b1111111111011111111111111111111111111111111111111111111111111111;
                endcase
            end
        endcase
    end
endmodule