
/**
 * @file class_hvec_gen_hdl.hpp
 * @brief This script generates HDL code for generating high-dimensional class vectors.
 * It is a novel method; for more information, please refer to our paper.
 *
 * @author Saeid Jamili and Marco Angioli
 * @note Author names are listed in alphabetical order.
 * @email <saeid.jamili@uniroma1.it>
 * @email <marco.angioli@uniroma1.it>
 *
 * @contributors
 *
 * @date Created: 24th July 2023
 * @date Last Updated: 23th August 2023
 *
 * @version 1.0.0
 *
 * @institute Sapienza University of Rome
 * @cite https://doi.org/10.xxxx/yyyyy
 *
 * @section DEPENDENCIES
 * - Dependency1: Description or version details.
 * - Dependency2: Description or version details.
 *
 * @section LICENSE
 * This file is part of the Aeneas HyperCompute Platform.
 *
 * Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 *
 * @section CHANGELOG
 * @version 1.0.0-dev - 23th August 2023
 * - Initial release
 *
 * @todo
 * - Complete level vector generator function
 * - Add training
 *
 * @see
 * -
 * -
 * -
 *
 */

module class_hvec_gen #(parameter int DI_PARALLEL_W_BITS = 64) (
  input logic [2:0] frame_id,
  input logic [1:0] frame_index,
  output logic [DI_PARALLEL_W_BITS-1:0] class_vec_out
);
  always_comb begin
    case (frame_id)
      0:
        case (frame_index)
          0:
            class_vec_out = 64'b010290861124500012451245952012451245084109939923124511310051106212210061512452360121701218124510161133572124501245124512151245124512450101245729690119510993124531825051412451245;
          1:
            class_vec_out = 64'b0208021122300022322221402232200402213210223208006019222200362233102090211223218213165223022322321322322322300223532150577018222361020111223223;
          2:
            class_vec_out = 64'b08505512600012612560012611803126120126690029119116006812637011501261268466110126012612612512612612605126138706490411261320058126126;
        endcase
      1:
        case (frame_index)
          0:
            class_vec_out = 64'b11501245123104135670200124512450124512101004551049614124510371245012454442124211094230124500117251612451228124518918124200124555100001212124501245124508471162064810071245124512451111;
          1:
            class_vec_out = 64'b159223223014118176002232230223221000161231372232092230223392221218530223002221012232112238822223002232270020122302232230172180079214223223223199;
          2:
            class_vec_out = 64'b91126113066431110012612601261260002111355126701260126068126110860126001155312611012654211260012628290011012601261260531180669412612612662;
        endcase
      2:
        case (frame_index)
          0:
            class_vec_out = 64'b0124512154100205123607812031012450123248598124501245123612451245102591796400077312451245028601099038511220012450124511751245823124524112341060158106312454784265124510405641245;
          1:
            class_vec_out = 64'b022321823001292220015509022302202189223022322022322313120112600035223223014021001692140022302231642234022394222901221972237202022314039223;
          2:
            class_vec_out = 64'b0126123190045124021030751260126333812601261001261267011810500093126126035011708999001260126951265712678108505811912696147712647060126;
        endcase
      3:
        case (frame_index)
          0:
            class_vec_out = 64'b012451238055812451239974012454288141229124550466709591245001245124512450122401245124512455291245124539212452412450100001730012451089124576112459746193011100172659124505463981245001150;
          1:
            class_vec_out = 64'b0223207094223221186022312019321822313014901552230022322322302210223223223572232234022332230218096102172112235222331925301340756622301102322300181;
          2:
            class_vec_out = 64'b0126123058126125790126651189812672990501260012612612601180126126126441261263512661260830620011895126691261584240116027511260227112600108;
        endcase
      4:
        case (frame_index)
          0:
            class_vec_out = 64'b063612450124510911730012450946124312119612450124536512450679501190124579401245103124501245124301245124512451053413348114531245124512450012451901245733136145146124512450124512450012451245;
          1:
            class_vec_out = 64'b027223022301990022309421125882230223302235144101802231280223922302232220223223223205511718602232232230022311822311407153223223022322300223223;
          2:
            class_vec_out = 64'b081126012611070012606812659401260126261265571301051268001264126012612501261241266462171061412612612600126331268010131126126012612600126126;
        endcase
      5:
        case (frame_index)
          0:
            class_vec_out = 64'b530904529167124535103358124512451245124505112205171245265120501118124584907250124512458820124501245745124512451196124500124500603100112431245951019357312451245123800071100153;
          1:
            class_vec_out = 64'b911294227223400257022322322322301921211022355222018822370033022322394022302234122322321222300223001811016522231210111032232232200101990069;
          2:
            class_vec_out = 64'b1411040211262402333126126126126071192912658990931267504801261261110126012682126126118126001260010416011201269805764126126126000680054;
        endcase
      6:
        case (frame_index)
          0:
            class_vec_out = 64'b61090007951245152003810481035124551245124502250123506684412451178012451245124571712251042354010880124512440012450394124511401245000119415354950108270122612450104101239;
          1:
            class_vec_out = 64'b51620063223720030219217223022322301090223032138223211022322322356218214146018502232210022301622310602230002236112107066021922302110223;
          2:
            class_vec_out = 64'b0113006912616008949712621261260640126029112664012612612693120781060890126118001260313126390126000116224452163101241260940119;
        endcase
      7:
        case (frame_index)
          0:
            class_vec_out = 64'b9418832381711245012457270124512320106811700012455101245124512455621245124512450605123629501244801245001219220115712451245106124512453462000124513124512450124512456391245421621000633;
          1:
            class_vec_out = 64'b21519055322302231150223222017020100223109223223223120223223223061223120022379223002183020522322342232236130002233223223022322318422316490000186;
          2:
            class_vec_out = 64'b97713820126012681012612601001080012655126126126102126126126032119190124481260010040122126126241261269440001264126126012612670126537830086;
        endcase
    endcase
  end
endmodule