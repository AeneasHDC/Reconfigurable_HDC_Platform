----
 -- @file level_hvec_gen_hdl.hpp
 -- @brief This script generates HDL code for generating high-dimensional LEVEL vectors.
 -- It is a novel method; for more information, please refer to our paper.
 --
 -- @author Saeid Jamili and Marco Angioli
 -- @note Author names are listed in alphabetical order.
 -- @email <saeid.jamili@uniroma1.it>
 -- @email <marco.angioli@uniroma1.it>
 --
 -- @contributors
 --
 -- @date Created: 24th July 2023
 -- @date Last Updated: 23th August 2023
 --
 -- @version 1.0.0
 --
 -- @institute Sapienza University of Rome
 -- @cite https://doi.org/10.xxxx/yyyyy
 --
 -- @section DEPENDENCIES
 -- - Dependency1: Description or version details.
 -- - Dependency2: Description or version details.
 --
 -- @section LICENSE
 -- This file is part of the Aeneas HyperCompute Platform.
 --
 -- Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 --
 -- @section CHANGELOG
 -- @version 1.0.0-dev - 23th August 2023
 -- - Initial release
 --
 -- @todo
 -- - Complete level vector generator function
 -- - Add training
 --
 -- @see
 -- -
 -- -
 -- -
 --
 --

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity level_vec_gen is
    Port ( level_vec_out : out  STD_LOGIC_VECTOR (63 downto 0);
           frame_index : in  STD_LOGIC_VECTOR (2 downto 0);
           frame_id : in  STD_LOGIC_VECTOR (4 downto 0));
end level_vec_gen;

architecture Behavioral of level_vec_gen is
begin
    process (frame_index, frame_id)
    begin
        -- Update this function to match your requirements
        case frame_index is
            when "000" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1000110001000110010100111010011110011001100111101100001011111001";
                    when "00001" => level_vec_out <= "1000110001000110010100111010011110011001100111101100001011111001";
                    when "00010" => level_vec_out <= "1000110001000110010100111010011110011001100111101100001011111001";
                    when "00011" => level_vec_out <= "1000110001000110010100111010011110011001100111101100001011111001";
                    when "00100" => level_vec_out <= "1000110001000110010100111011011110011001100111101100001011111001";
                    when "00101" => level_vec_out <= "1000110001010110010100111011011110011101100111101100001011111001";
                    when "00110" => level_vec_out <= "1000110001010110010100111011011110011101100111101100011011111001";
                    when "00111" => level_vec_out <= "1000110001010110010100111011011110111101100111101100011011111011";
                    when "01000" => level_vec_out <= "1000110101010110010100111011011110111101100111101100011011111011";
                    when "01001" => level_vec_out <= "1000110101010110010100111011011110111101100111101100011011111011";
                    when "01010" => level_vec_out <= "1000110101010110010100111011011110111101100111101100011011111011";
                    when "01011" => level_vec_out <= "1000110101010110010100111011011110111101100111101100011011111011";
                    when "01100" => level_vec_out <= "1000110101010110011100111011011110111101110111101110011011111111";
                    when "01101" => level_vec_out <= "1000110101011110011100111011011110111101110111101110011011111111";
                    when "01110" => level_vec_out <= "1000110101011110011100111011011110111101110111101110011011111111";
                    when "01111" => level_vec_out <= "1000110101011110011100111011011110111101110111101110011011111111";
                    when "10000" => level_vec_out <= "1100110101011110011100111011011110111101110111111110011011111111";
                    when "10001" => level_vec_out <= "1100110101011110011100111011011111111101110111111110011011111111";
                    when "10010" => level_vec_out <= "1100110101011111011100111011011111111111110111111110011011111111";
                    when "10011" => level_vec_out <= "1100110101011111011100111011011111111111110111111111011011111111";
                    when "10100" => level_vec_out <= "1100110101111111011100111011011111111111110111111111011011111111";
                    when "10101" => level_vec_out <= "1100110101111111011100111011011111111111110111111111011011111111";
                    when "10110" => level_vec_out <= "1100110101111111011101111111011111111111110111111111111011111111";
                    when "10111" => level_vec_out <= "1100110101111111011101111111011111111111111111111111111011111111";
                    when "11000" => level_vec_out <= "1100110101111111011101111111011111111111111111111111111011111111";
                    when "11001" => level_vec_out <= "1100110101111111111101111111011111111111111111111111111111111111";
                    when "11010" => level_vec_out <= "1100111101111111111101111111011111111111111111111111111111111111";
                    when "11011" => level_vec_out <= "1100111101111111111101111111111111111111111111111111111111111111";
                    when "11100" => level_vec_out <= "1100111111111111111101111111111111111111111111111111111111111111";
                    when "11101" => level_vec_out <= "1100111111111111111101111111111111111111111111111111111111111111";
                    when "11110" => level_vec_out <= "1101111111111111111111111111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "001" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1010001010001000110101011111110010110010101001111010110111010101";
                    when "00001" => level_vec_out <= "1010001010001001110101011111111010110010101001111010110111010101";
                    when "00010" => level_vec_out <= "1010001010001001110101011111111010110010101001111010111111010101";
                    when "00011" => level_vec_out <= "1010001010001001110101011111111010110010101001111010111111010101";
                    when "00100" => level_vec_out <= "1010001010001001110101011111111010110010111001111010111111010111";
                    when "00101" => level_vec_out <= "1010001010001001110101011111111010110010111001111010111111010111";
                    when "00110" => level_vec_out <= "1010001010001001110101011111111010110010111001111010111111010111";
                    when "00111" => level_vec_out <= "1010001010011001110101011111111010110010111001111010111111010111";
                    when "01000" => level_vec_out <= "1010001010011001110101011111111010110010111001111010111111010111";
                    when "01001" => level_vec_out <= "1010011010011001110101011111111010110010111001111010111111010111";
                    when "01010" => level_vec_out <= "1010011010011001110101011111111010110010111001111010111111110111";
                    when "01011" => level_vec_out <= "1010011010011001110101011111111010110010111001111010111111110111";
                    when "01100" => level_vec_out <= "1010011011011001110101011111111010110010111001111010111111110111";
                    when "01101" => level_vec_out <= "1110011011011001110101011111111010110010111001111011111111110111";
                    when "01110" => level_vec_out <= "1110011011011001110101011111111010110010111001111011111111110111";
                    when "01111" => level_vec_out <= "1110111011011001111101011111111010110010111001111011111111111111";
                    when "10000" => level_vec_out <= "1110111111011001111101011111111010110110111001111011111111111111";
                    when "10001" => level_vec_out <= "1110111111011001111101011111111010110110111001111011111111111111";
                    when "10010" => level_vec_out <= "1110111111011001111101011111111010110110111001111011111111111111";
                    when "10011" => level_vec_out <= "1110111111011001111101011111111010110110111001111011111111111111";
                    when "10100" => level_vec_out <= "1111111111011001111101011111111010110110111001111011111111111111";
                    when "10101" => level_vec_out <= "1111111111111001111101011111111110110110111001111011111111111111";
                    when "10110" => level_vec_out <= "1111111111111001111101011111111111110110111101111011111111111111";
                    when "10111" => level_vec_out <= "1111111111111001111101011111111111110110111101111011111111111111";
                    when "11000" => level_vec_out <= "1111111111111001111101111111111111110110111111111011111111111111";
                    when "11001" => level_vec_out <= "1111111111111001111101111111111111111110111111111011111111111111";
                    when "11010" => level_vec_out <= "1111111111111001111101111111111111111110111111111011111111111111";
                    when "11011" => level_vec_out <= "1111111111111001111101111111111111111110111111111011111111111111";
                    when "11100" => level_vec_out <= "1111111111111001111111111111111111111111111111111011111111111111";
                    when "11101" => level_vec_out <= "1111111111111001111111111111111111111111111111111111111111111111";
                    when "11110" => level_vec_out <= "1111111111111001111111111111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111011111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "010" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0111001110010010101110110001111011011101111011011111100001111011";
                    when "00001" => level_vec_out <= "1111001110010010101110110001111011011101111011011111100001111011";
                    when "00010" => level_vec_out <= "1111001110010010101110110001111011011101111011011111100101111011";
                    when "00011" => level_vec_out <= "1111001110010010101110110001111011011101111111011111100101111011";
                    when "00100" => level_vec_out <= "1111001110010010101110110001111011011101111111011111100101111011";
                    when "00101" => level_vec_out <= "1111001110010010101110110001111011011111111111011111100101111011";
                    when "00110" => level_vec_out <= "1111001110010010101110110001111011011111111111011111100101111011";
                    when "00111" => level_vec_out <= "1111001110010010101110110001111011011111111111011111100101111011";
                    when "01000" => level_vec_out <= "1111001110110010101110110011111011011111111111011111100101111011";
                    when "01001" => level_vec_out <= "1111001110110010101110110011111011011111111111011111110101111011";
                    when "01010" => level_vec_out <= "1111001110110010111110111011111011011111111111011111111101111011";
                    when "01011" => level_vec_out <= "1111001110110010111110111011111011111111111111011111111101111011";
                    when "01100" => level_vec_out <= "1111001110110010111110111011111011111111111111011111111101111011";
                    when "01101" => level_vec_out <= "1111001110110010111110111011111011111111111111011111111101111011";
                    when "01110" => level_vec_out <= "1111001110110010111110111011111011111111111111011111111101111011";
                    when "01111" => level_vec_out <= "1111001110110010111110111011111011111111111111011111111101111011";
                    when "10000" => level_vec_out <= "1111001110110010111110111011111011111111111111011111111101111011";
                    when "10001" => level_vec_out <= "1111001110110010111111111011111011111111111111011111111101111011";
                    when "10010" => level_vec_out <= "1111001110110010111111111011111011111111111111011111111101111011";
                    when "10011" => level_vec_out <= "1111001110110010111111111011111011111111111111011111111101111011";
                    when "10100" => level_vec_out <= "1111001110110010111111111011111011111111111111011111111101111111";
                    when "10101" => level_vec_out <= "1111001110110011111111111011111011111111111111111111111101111111";
                    when "10110" => level_vec_out <= "1111001110110011111111111011111011111111111111111111111101111111";
                    when "10111" => level_vec_out <= "1111001110110011111111111011111111111111111111111111111101111111";
                    when "11000" => level_vec_out <= "1111001111110111111111111011111111111111111111111111111101111111";
                    when "11001" => level_vec_out <= "1111101111111111111111111011111111111111111111111111111101111111";
                    when "11010" => level_vec_out <= "1111101111111111111111111011111111111111111111111111111101111111";
                    when "11011" => level_vec_out <= "1111101111111111111111111011111111111111111111111111111101111111";
                    when "11100" => level_vec_out <= "1111101111111111111111111111111111111111111111111111111101111111";
                    when "11101" => level_vec_out <= "1111101111111111111111111111111111111111111111111111111101111111";
                    when "11110" => level_vec_out <= "1111101111111111111111111111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "011" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0111111001001100111101100100000010111010000100011001011100011001";
                    when "00001" => level_vec_out <= "0111111001001100111101100100000010111010000100011001011100011001";
                    when "00010" => level_vec_out <= "0111111001001100111101100100000010111010010100011001011100011001";
                    when "00011" => level_vec_out <= "0111111001101100111101100100000010111010111100011001011100011101";
                    when "00100" => level_vec_out <= "0111111001101100111101100100000010111010111100011001011110011101";
                    when "00101" => level_vec_out <= "0111111001101100111101100100000010111010111100011001111110011101";
                    when "00110" => level_vec_out <= "0111111011101100111101101100000010111010111100011001111111011101";
                    when "00111" => level_vec_out <= "0111111011101100111101101100000010111010111100011001111111111101";
                    when "01000" => level_vec_out <= "0111111011101100111101101100000010111010111110111001111111111101";
                    when "01001" => level_vec_out <= "0111111011101100111101101110000010111010111110111001111111111101";
                    when "01010" => level_vec_out <= "0111111011101100111101101110000010111010111110111001111111111101";
                    when "01011" => level_vec_out <= "0111111011101100111101101110000010111010111110111001111111111101";
                    when "01100" => level_vec_out <= "0111111011101100111101101110000010111010111110111011111111111101";
                    when "01101" => level_vec_out <= "0111111011101100111101101110000010111010111110111011111111111101";
                    when "01110" => level_vec_out <= "0111111011101100111101101110100010111010111110111011111111111101";
                    when "01111" => level_vec_out <= "0111111011101100111101101110100010111010111110111011111111111101";
                    when "10000" => level_vec_out <= "0111111011101100111101101110100010111010111110111011111111111101";
                    when "10001" => level_vec_out <= "0111111111101100111111101110100010111010111110111011111111111101";
                    when "10010" => level_vec_out <= "0111111111111100111111101110100110111010111111111011111111111101";
                    when "10011" => level_vec_out <= "0111111111111110111111101110100110111010111111111011111111111101";
                    when "10100" => level_vec_out <= "0111111111111110111111101110100110111010111111111011111111111101";
                    when "10101" => level_vec_out <= "0111111111111110111111101110100110111110111111111011111111111101";
                    when "10110" => level_vec_out <= "0111111111111110111111101110100110111110111111111011111111111111";
                    when "10111" => level_vec_out <= "1111111111111110111111101110100110111110111111111011111111111111";
                    when "11000" => level_vec_out <= "1111111111111110111111101110101110111110111111111011111111111111";
                    when "11001" => level_vec_out <= "1111111111111110111111101110101110111110111111111011111111111111";
                    when "11010" => level_vec_out <= "1111111111111110111111101110101110111110111111111111111111111111";
                    when "11011" => level_vec_out <= "1111111111111110111111101110101110111110111111111111111111111111";
                    when "11100" => level_vec_out <= "1111111111111111111111111110101110111110111111111111111111111111";
                    when "11101" => level_vec_out <= "1111111111111111111111111110101111111110111111111111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111110101111111110111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111110101111111111111111111111111111111111";
                when others => null;
                end case;
            when "100" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0101000001111110110001011000111001010111110010010001100100101000";
                    when "00001" => level_vec_out <= "0101000001111110110101011010111001010111110010011001100100101000";
                    when "00010" => level_vec_out <= "0101000001111110110101011010111001010111110010011001100100101001";
                    when "00011" => level_vec_out <= "0101000001111110110101011010111001010111111010011001100100101001";
                    when "00100" => level_vec_out <= "0101000001111110110101011010111001010111111111011001100100101001";
                    when "00101" => level_vec_out <= "0101000001111110110101011011111011010111111111011001100100101001";
                    when "00110" => level_vec_out <= "0101000001111110110101011011111011010111111111011001100100101001";
                    when "00111" => level_vec_out <= "0101000001111110110101011011111011010111111111111001100100101001";
                    when "01000" => level_vec_out <= "0101000001111110110101011011111011010111111111111001100100101001";
                    when "01001" => level_vec_out <= "0101000001111110110101011011111011010111111111111001110100101001";
                    when "01010" => level_vec_out <= "0101000001111110110101011011111111010111111111111001110100101011";
                    when "01011" => level_vec_out <= "0101000001111110110101011011111111010111111111111011110100101011";
                    when "01100" => level_vec_out <= "0101000001111110110101011011111111010111111111111011110100101011";
                    when "01101" => level_vec_out <= "0101000001111110110101011011111111010111111111111011110110101011";
                    when "01110" => level_vec_out <= "0101010001111110110111011011111111011111111111111011110110101011";
                    when "01111" => level_vec_out <= "0101010001111110110111011111111111011111111111111011110110101011";
                    when "10000" => level_vec_out <= "0101010101111110110111011111111111011111111111111011110110101011";
                    when "10001" => level_vec_out <= "0101010101111110110111011111111111111111111111111011110110111011";
                    when "10010" => level_vec_out <= "0101010101111110110111011111111111111111111111111011110110111011";
                    when "10011" => level_vec_out <= "0101010101111110110111011111111111111111111111111011111110111011";
                    when "10100" => level_vec_out <= "0101010101111110110111011111111111111111111111111011111110111011";
                    when "10101" => level_vec_out <= "0101010101111110110111011111111111111111111111111011111110111011";
                    when "10110" => level_vec_out <= "0101010101111110110111011111111111111111111111111011111110111111";
                    when "10111" => level_vec_out <= "0101011101111110110111011111111111111111111111111011111110111111";
                    when "11000" => level_vec_out <= "0101011101111110110111011111111111111111111111111011111110111111";
                    when "11001" => level_vec_out <= "0101011101111110110111011111111111111111111111111011111110111111";
                    when "11010" => level_vec_out <= "0101011101111111110111011111111111111111111111111011111110111111";
                    when "11011" => level_vec_out <= "1111011101111111111111111111111111111111111111111011111110111111";
                    when "11100" => level_vec_out <= "1111111101111111111111111111111111111111111111111011111110111111";
                    when "11101" => level_vec_out <= "1111111101111111111111111111111111111111111111111011111110111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111110111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111110111111";
                when others => null;
                end case;
            when "101" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1101100000010001101011001001110101000111010001100110101110010010";
                    when "00001" => level_vec_out <= "1101100000010001101011001001110101000111010001100110101110010010";
                    when "00010" => level_vec_out <= "1101100000010011101011101001111101000111010001100110101110010010";
                    when "00011" => level_vec_out <= "1101100000010011101011101001111101000111010001110110101110010010";
                    when "00100" => level_vec_out <= "1101100000010011101011101001111101000111010001110110101110010010";
                    when "00101" => level_vec_out <= "1101100000010011101011101001111101000111010001110110101110010010";
                    when "00110" => level_vec_out <= "1101100000010011101011101001111101000111010001110111101110010010";
                    when "00111" => level_vec_out <= "1101100000010111101011101001111101000111010001110111101110010010";
                    when "01000" => level_vec_out <= "1101100000010111101011101001111101000111010001110111111110010010";
                    when "01001" => level_vec_out <= "1101100000010111101011101001111101000111010001110111111110010011";
                    when "01010" => level_vec_out <= "1101100000010111101011101001111101000111010001110111111110010011";
                    when "01011" => level_vec_out <= "1101100000010111101011101001111101000111110001111111111110010011";
                    when "01100" => level_vec_out <= "1101100000010111101011101001111101000111110001111111111110010111";
                    when "01101" => level_vec_out <= "1101100000011111101011101001111101000111111001111111111110010111";
                    when "01110" => level_vec_out <= "1101110000011111101111101001111101010111111001111111111110010111";
                    when "01111" => level_vec_out <= "1101110100011111101111101001111101011111111001111111111110010111";
                    when "10000" => level_vec_out <= "1101110100011111101111101001111101011111111001111111111110110111";
                    when "10001" => level_vec_out <= "1101110100011111101111101001111101011111111001111111111110110111";
                    when "10010" => level_vec_out <= "1101110100011111101111101001111101011111111001111111111110110111";
                    when "10011" => level_vec_out <= "1101110100011111101111101001111101111111111001111111111111110111";
                    when "10100" => level_vec_out <= "1101110100011111101111101001111101111111111001111111111111110111";
                    when "10101" => level_vec_out <= "1101110100011111101111101001111101111111111001111111111111110111";
                    when "10110" => level_vec_out <= "1101110100011111101111101001111101111111111001111111111111110111";
                    when "10111" => level_vec_out <= "1101110110011111101111101001111101111111111001111111111111110111";
                    when "11000" => level_vec_out <= "1101110110011111101111101101111111111111111011111111111111110111";
                    when "11001" => level_vec_out <= "1101110110111111111111101101111111111111111011111111111111110111";
                    when "11010" => level_vec_out <= "1101110111111111111111101101111111111111111011111111111111110111";
                    when "11011" => level_vec_out <= "1111110111111111111111101101111111111111111011111111111111110111";
                    when "11100" => level_vec_out <= "1111110111111111111111111101111111111111111011111111111111110111";
                    when "11101" => level_vec_out <= "1111111111111111111111111101111111111111111011111111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111111011111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111011111111111111111111";
                when others => null;
                end case;
            when "110" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0100010101100101110000010010011010011000100100111110101100001111";
                    when "00001" => level_vec_out <= "0100010101100101110000010010011010011000101100111110101100001111";
                    when "00010" => level_vec_out <= "0100010101100101110000010010011010011000101101111110101100001111";
                    when "00011" => level_vec_out <= "0100010101110101110000010010011010011000101101111110101100001111";
                    when "00100" => level_vec_out <= "0100011101110101110000110010011010011000101101111110101100001111";
                    when "00101" => level_vec_out <= "0100011101110101110000110010011010011000101101111110101100001111";
                    when "00110" => level_vec_out <= "0100011101110101110000110010011010011000101101111110101100001111";
                    when "00111" => level_vec_out <= "0100011101110101110010110010011010011000101101111110101100101111";
                    when "01000" => level_vec_out <= "0100011101110101110010110010011011011000101101111110101100101111";
                    when "01001" => level_vec_out <= "0100011101110101110010110110011011011000101101111110101100101111";
                    when "01010" => level_vec_out <= "0100011101110101110010110111011011011000101101111110101110101111";
                    when "01011" => level_vec_out <= "0100011111110101110011110111011011011000101101111110101110101111";
                    when "01100" => level_vec_out <= "0100011111110101110011110111011011011000101101111110101110101111";
                    when "01101" => level_vec_out <= "0100011111110101110011110111011011011000101101111110101110101111";
                    when "01110" => level_vec_out <= "0100011111110101110011110111011011011000101101111110101110101111";
                    when "01111" => level_vec_out <= "0100011111110101110011110111011011011000101101111110101110101111";
                    when "10000" => level_vec_out <= "0100011111110101110011110111011011011000101101111110101111101111";
                    when "10001" => level_vec_out <= "0100011111110111110011110111011011011000101101111110101111101111";
                    when "10010" => level_vec_out <= "0100011111110111110111110111011011011000101101111110101111101111";
                    when "10011" => level_vec_out <= "0100011111110111110111110111011011011000101111111110101111101111";
                    when "10100" => level_vec_out <= "0100011111110111110111111111011111011000101111111111101111111111";
                    when "10101" => level_vec_out <= "0100011111110111110111111111011111011000101111111111101111111111";
                    when "10110" => level_vec_out <= "0100011111110111110111111111011111011000101111111111101111111111";
                    when "10111" => level_vec_out <= "0110011111111111110111111111011111011000101111111111101111111111";
                    when "11000" => level_vec_out <= "0110011111111111110111111111011111011000101111111111101111111111";
                    when "11001" => level_vec_out <= "0110011111111111110111111111011111011010101111111111101111111111";
                    when "11010" => level_vec_out <= "0110011111111111111111111111011111111010111111111111111111111111";
                    when "11011" => level_vec_out <= "0110011111111111111111111111011111111011111111111111111111111111";
                    when "11100" => level_vec_out <= "0110011111111111111111111111011111111011111111111111111111111111";
                    when "11101" => level_vec_out <= "1110011111111111111111111111011111111011111111111111111111111111";
                    when "11110" => level_vec_out <= "1110011111111111111111111111011111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111011111111111111111111111111111111111";
                when others => null;
                end case;
            when "111" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0100000110000011111000100000110010001010100000011000111011110101";
                    when "00001" => level_vec_out <= "0100000110000011111000100000110010001010100010011000111011110101";
                    when "00010" => level_vec_out <= "0100000110000011111000100000110010001010100010011000111011110101";
                    when "00011" => level_vec_out <= "0100000110000011111000100000110010001010100010011000111011110101";
                    when "00100" => level_vec_out <= "0100000110000011111000100000110010001010100010011000111011110101";
                    when "00101" => level_vec_out <= "0100000110000011111001100000110010001010100010011000111011110111";
                    when "00110" => level_vec_out <= "0100000110000011111001101000111010001010100011011000111011110111";
                    when "00111" => level_vec_out <= "0100000110000011111001101000111010001010100011011000111011110111";
                    when "01000" => level_vec_out <= "0100000110010011111001101000111010001010100011011000111011110111";
                    when "01001" => level_vec_out <= "0100000110010011111001101000111010001010100111011000111011111111";
                    when "01010" => level_vec_out <= "0100000110010011111001101000111010001010100111011000111011111111";
                    when "01011" => level_vec_out <= "0101000110010011111001101000111010001010100111011000111111111111";
                    when "01100" => level_vec_out <= "0101000110010011111001101000111010101010100111011000111111111111";
                    when "01101" => level_vec_out <= "0101000110010011111101101000111010101010100111111000111111111111";
                    when "01110" => level_vec_out <= "0101000110010011111101101000111010101110100111111000111111111111";
                    when "01111" => level_vec_out <= "1101000110010011111101111000111010101110100111111000111111111111";
                    when "10000" => level_vec_out <= "1101000110010011111101111000111010101111100111111000111111111111";
                    when "10001" => level_vec_out <= "1101000110010011111101111000111010111111100111111000111111111111";
                    when "10010" => level_vec_out <= "1101000110010011111101111000111010111111110111111100111111111111";
                    when "10011" => level_vec_out <= "1101000110010111111101111010111010111111110111111100111111111111";
                    when "10100" => level_vec_out <= "1101000110011111111101111010111010111111110111111100111111111111";
                    when "10101" => level_vec_out <= "1101000111011111111101111010111010111111111111111101111111111111";
                    when "10110" => level_vec_out <= "1101000111011111111101111010111110111111111111111101111111111111";
                    when "10111" => level_vec_out <= "1101010111011111111101111010111110111111111111111101111111111111";
                    when "11000" => level_vec_out <= "1101010111011111111101111010111110111111111111111101111111111111";
                    when "11001" => level_vec_out <= "1101010111011111111101111010111110111111111111111101111111111111";
                    when "11010" => level_vec_out <= "1101010111011111111101111010111110111111111111111101111111111111";
                    when "11011" => level_vec_out <= "1101010111011111111101111010111110111111111111111111111111111111";
                    when "11100" => level_vec_out <= "1101010111011111111101111010111110111111111111111111111111111111";
                    when "11101" => level_vec_out <= "1111110111011111111101111110111110111111111111111111111111111111";
                    when "11110" => level_vec_out <= "1111110111011111111111111110111110111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111110111011111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when others => null;
        end case;
    end process;
end Behavioral;