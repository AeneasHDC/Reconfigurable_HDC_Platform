/**
 * @file level_hvec_gen_hdl.hpp
 * @brief This script generates HDL code for generating high-dimensional LEVEL vectors.
 * It is a novel method; for more information, please refer to our paper.
 *
 * @author Saeid Jamili and Marco Angioli
 * @note Author names are listed in alphabetical order.
 * @email <saeid.jamili@uniroma1.it>
 * @email <marco.angioli@uniroma1.it>
 *
 * @contributors
 *
 * @date Created: 24th July 2023
 * @date Last Updated: 23th August 2023
 *
 * @version 0.0.1-dev
 *
 * @institute Sapienza University of Rome
 * @cite https://doi.org/10.xxxx/yyyyy
 *
 * @section DEPENDENCIES
 * - Dependency1: Description or version details.
 * - Dependency2: Description or version details.
 *
 * @section LICENSE
 * This file is part of the Aeneas HyperCompute Platform.
 *
 * Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 *
 * @section CHANGELOG
 * @version 1.0.0-dev - 23th August 2023
 * - Initial release
 *
 * @todo
 * - Complete level vector generator function
 * - Add training
 *
 * @see
 * -
 * -
 * -
 *
 */

module level_vec_gen (
    output reg [99:0] level_vec_out,
    input [3:0] frame_index,
    input [4:0] frame_id
);
    always @(*) begin
        // Update this function to match your requirements
        case (frame_index)
            0: begin
                case (frame_id)
                    0: level_vec_out = 100'b0011100101100010100111001000010110101110010001010000100101110011010001011110011001010001100000111110;
                    1: level_vec_out = 100'b0011100101100010100111001000010110101110010001010000100101110011011001011110011011010001100000111110;
                    2: level_vec_out = 100'b0011100101100010100111001000010110101110010001010000100101110011011001011111011011011001100000111110;
                    3: level_vec_out = 100'b0011100101100010100111001000010110101110010001010000100101110011111001011111011011011001100000111110;
                    4: level_vec_out = 100'b0011100101100010100111001000010110101110010001010000100101110011111001011111011011011001100010111111;
                    5: level_vec_out = 100'b0011100101100010100111001100010110101110010001010000100101110011111001011111011011111001100010111111;
                    6: level_vec_out = 100'b0011110101100010100111001100010110101110010001010000100101110011111001011111011011111101100010111111;
                    7: level_vec_out = 100'b0011110101100010100111001100010110101110010001110000100101110011111001011111011011111101100010111111;
                    8: level_vec_out = 100'b0011110101100010100111001100010110101110110001110000100101110011111001011111011011111101100010111111;
                    9: level_vec_out = 100'b1011110101100010100111001100010110101110110001110000100101110011111001011111011011111101101010111111;
                    10: level_vec_out = 100'b1011110101100010100111001100010110101110110001110010100101110011111001011111011011111101101010111111;
                    11: level_vec_out = 100'b1011110101100010100111101100110110101110110011110010100101110011111001011111011011111101101010111111;
                    12: level_vec_out = 100'b1011110101100010100111101100110110101110110011110010100101110111111101011111011011111101101010111111;
                    13: level_vec_out = 100'b1011110101101010100111101100110110101110110011110010100101110111111101011111011111111101101011111111;
                    14: level_vec_out = 100'b1011110101101010101111101100110110101111110011110010100101110111111101011111011111111101101011111111;
                    15: level_vec_out = 100'b1011110101101010101111101100110110101111110011111010100101110111111101011111111111111101101011111111;
                    16: level_vec_out = 100'b1011110101111010101111101100110110101111110011111010100101111111111101011111111111111101101011111111;
                    17: level_vec_out = 100'b1011111101111010101111101100110110101111110011111010100101111111111101011111111111111101101011111111;
                    18: level_vec_out = 100'b1011111111111010101111101100110110101111110011111010110101111111111101011111111111111101101011111111;
                    19: level_vec_out = 100'b1011111111111010101111101100110110101111111011111010111101111111111111011111111111111101101011111111;
                    20: level_vec_out = 100'b1011111111111010101111101110110110101111111011111010111101111111111111011111111111111101101011111111;
                    21: level_vec_out = 100'b1011111111111010101111101110110110101111111011111010111101111111111111011111111111111101101011111111;
                    22: level_vec_out = 100'b1011111111111010101111101110110110101111111011111010111111111111111111011111111111111101101011111111;
                    23: level_vec_out = 100'b1011111111111010111111101110110110101111111111111010111111111111111111011111111111111101101011111111;
                    24: level_vec_out = 100'b1011111111111010111111101110111110101111111111111010111111111111111111011111111111111101101111111111;
                    25: level_vec_out = 100'b1011111111111110111111101110111110101111111111111010111111111111111111111111111111111101101111111111;
                    26: level_vec_out = 100'b1011111111111110111111101110111110101111111111111011111111111111111111111111111111111101101111111111;
                    27: level_vec_out = 100'b1011111111111110111111101110111111101111111111111011111111111111111111111111111111111101111111111111;
                    28: level_vec_out = 100'b1111111111111110111111101110111111101111111111111111111111111111111111111111111111111111111111111111;
                    29: level_vec_out = 100'b1111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111;
                endcase
            end
            1: begin
                case (frame_id)
                    0: level_vec_out = 100'b1000011000010101010110001011010100010000100101100110111110001101111100101110101111001110011111101100;
                    1: level_vec_out = 100'b1100011001010101010110001011010100010000100101100110111110001101111100101110101111001110011111101100;
                    2: level_vec_out = 100'b1100011001010101010110101011010100010000100111100110111110001101111100101110101111001110011111101100;
                    3: level_vec_out = 100'b1100011001010101010110101011010100010000100111100110111110001101111100101110101111011111011111101100;
                    4: level_vec_out = 100'b1101011001010101010110101011010100010000100111100110111110101101111100101110101111011111011111101100;
                    5: level_vec_out = 100'b1101111001010101010110101011011100010000100111100110111110101101111100101110101111011111011111101100;
                    6: level_vec_out = 100'b1101111001010101010110101011011100010000100111100110111110101101111100101110101111011111011111101100;
                    7: level_vec_out = 100'b1101111001010101010111101011011100010000100111100110111110101101111100101110101111011111011111101100;
                    8: level_vec_out = 100'b1101111001010101010111101011011100010000100111100110111110101101111100101110101111011111111111101100;
                    9: level_vec_out = 100'b1101111011010101010111101011011100010000100111100110111110101101111100101110101111011111111111101100;
                    10: level_vec_out = 100'b1101111011010101010111101011011100010000100111100110111110101101111100101110101111011111111111101100;
                    11: level_vec_out = 100'b1101111011010101010111101011011100010000100111100110111110101101111100101110101111011111111111101100;
                    12: level_vec_out = 100'b1101111011010101010111101011011100010010100111100110111110101101111100101110101111011111111111101100;
                    13: level_vec_out = 100'b1101111011010101010111101011011100010010100111100110111110101101111100101110101111011111111111101100;
                    14: level_vec_out = 100'b1101111011011101010111101011011100010010100111100110111110101101111100101110101111111111111111101100;
                    15: level_vec_out = 100'b1101111011011101010111101011011100010010100111100110111110101101111100101110101111111111111111101100;
                    16: level_vec_out = 100'b1101111011011101010111101011011110010110100111100110111110101101111100101110101111111111111111101100;
                    17: level_vec_out = 100'b1101111011011101010111101011011110011110100111100110111110101101111100101110101111111111111111101100;
                    18: level_vec_out = 100'b1101111011011101011111101011011110011110100111100110111110101101111100101110101111111111111111101100;
                    19: level_vec_out = 100'b1101111011011101011111101011011110011110100111100110111111101101111100101110101111111111111111101100;
                    20: level_vec_out = 100'b1101111011011101011111101011111110011110100111100110111111101101111100101110101111111111111111101110;
                    21: level_vec_out = 100'b1101111011011101111111101011111110011110100111100110111111101101111100101110101111111111111111101110;
                    22: level_vec_out = 100'b1101111111111101111111101011111110011110100111100110111111101101111100101110101111111111111111101110;
                    23: level_vec_out = 100'b1101111111111111111111101111111110011110100111100111111111101101111110101110101111111111111111101110;
                    24: level_vec_out = 100'b1101111111111111111111101111111110011111100111100111111111101101111110101111101111111111111111101110;
                    25: level_vec_out = 100'b1111111111111111111111101111111110011111101111100111111111101101111110111111101111111111111111101111;
                    26: level_vec_out = 100'b1111111111111111111111101111111110011111101111110111111111101101111110111111101111111111111111101111;
                    27: level_vec_out = 100'b1111111111111111111111111111111110111111101111110111111111101101111110111111101111111111111111101111;
                    28: level_vec_out = 100'b1111111111111111111111111111111110111111101111110111111111101101111110111111101111111111111111111111;
                    29: level_vec_out = 100'b1111111111111111111111111111111111111111101111110111111111101101111111111111101111111111111111111111;
                endcase
            end
            2: begin
                case (frame_id)
                    0: level_vec_out = 100'b0100010100011101001000010001100111011001000110010111011000100010100111110111100110011001100111100011;
                    1: level_vec_out = 100'b0100010100011101001000010011100111011001000110010111011000100010100111110111100110011001100111100011;
                    2: level_vec_out = 100'b0100010100011101001000010011100111011001000110010111011100100010100111110111100110011001100111100011;
                    3: level_vec_out = 100'b0100010100011101001000010011100111011001000110010111011100100010100111110111100110011001100111100011;
                    4: level_vec_out = 100'b0100010100011101001000010011100111011001000110010111011100100010100111110111100110011001100111100011;
                    5: level_vec_out = 100'b0100010100011101001000010011100111011001000110110111011100100010100111110111100110011001100111101011;
                    6: level_vec_out = 100'b0100010110011101001000010011100111011001000111110111011100100010100111110111100110011101100111101011;
                    7: level_vec_out = 100'b0100010110011101001000110011100111011001000111110111011100100010100111110111100110011101100111101011;
                    8: level_vec_out = 100'b0100010110011101001000110011100111011001000111110111011100100010100111110111100110011101100111101011;
                    9: level_vec_out = 100'b0100010110011101001000110011100111011001000111110111011100100010100111110111100110011101100111101011;
                    10: level_vec_out = 100'b0100010110011101101000110011100111011001000111110111011100101010100111110111100110011101100111101011;
                    11: level_vec_out = 100'b0100110110011101101000110011110111011001000111110111011100101010100111110111100110011101100111101011;
                    12: level_vec_out = 100'b0100110110011101101000110011110111011001001111110111011100101010110111110111100111011101100111101111;
                    13: level_vec_out = 100'b0100110110011101101000110011110111011001001111110111011100101010110111110111100111011101100111101111;
                    14: level_vec_out = 100'b0100110110011101101000110011110111011001001111110111111100101010110111110111100111011101100111101111;
                    15: level_vec_out = 100'b0100110110011101101000110011110111011001001111110111111100101010110111110111100111011101100111101111;
                    16: level_vec_out = 100'b0100110110011101101000110011110111011001001111110111111100101010110111110111100111011101100111101111;
                    17: level_vec_out = 100'b0100110110011101101000110011110111111001001111110111111100101010110111110111110111011101100111101111;
                    18: level_vec_out = 100'b0101110110011101101000110011110111111001001111111111111110101110110111110111110111011111100111101111;
                    19: level_vec_out = 100'b1101111110011101101000110011111111111011001111111111111110101110110111110111111111011111100111101111;
                    20: level_vec_out = 100'b1101111110011101101000110011111111111011001111111111111110111110110111111111111111111111100111101111;
                    21: level_vec_out = 100'b1101111110011101101000110011111111111011001111111111111110111110111111111111111111111111100111101111;
                    22: level_vec_out = 100'b1101111110011101101000110011111111111011001111111111111110111110111111111111111111111111100111101111;
                    23: level_vec_out = 100'b1101111110011111101000110011111111111111001111111111111110111110111111111111111111111111100111101111;
                    24: level_vec_out = 100'b1101111110011111101000110011111111111111101111111111111110111110111111111111111111111111100111101111;
                    25: level_vec_out = 100'b1101111110011111101000110011111111111111111111111111111110111110111111111111111111111111101111101111;
                    26: level_vec_out = 100'b1101111110011111101101110011111111111111111111111111111111111110111111111111111111111111111111101111;
                    27: level_vec_out = 100'b1101111110011111101101111011111111111111111111111111111111111111111111111111111111111111111111101111;
                    28: level_vec_out = 100'b1101111110011111101101111011111111111111111111111111111111111111111111111111111111111111111111101111;
                    29: level_vec_out = 100'b1111111111011111101101111011111111111111111111111111111111111111111111111111111111111111111111101111;
                endcase
            end
            3: begin
                case (frame_id)
                    0: level_vec_out = 100'b1110100001011101100011001010011101101000100111100100010101101011111001101001111001101100010111100010;
                    1: level_vec_out = 100'b1110100001011101100011001010011101101000100111100100010101101011111001101001111001101100010111100010;
                    2: level_vec_out = 100'b1110100001011101100011001010011101101000100111100100010101101011111001101001111001101100010111100010;
                    3: level_vec_out = 100'b1110100001011101100011001010011101101000100111100100010101101011111001101001111001101101010111100110;
                    4: level_vec_out = 100'b1111101001011101100011001010011101101010100111100100010101101011111001101001111001101101010111100111;
                    5: level_vec_out = 100'b1111101001011101100011001010011101101010100111100100010101101011111001101001111001101101010111101111;
                    6: level_vec_out = 100'b1111101001111101100011001010011101101010100111100101010101101011111001101001111001101101011111101111;
                    7: level_vec_out = 100'b1111101001111101101011001010011101101010100111100101010101101011111001101101111001101101011111101111;
                    8: level_vec_out = 100'b1111111001111101101011001010011101101010100111100101010101101011111001101101111001101101011111101111;
                    9: level_vec_out = 100'b1111111001111101101011001010111101101010100111100101010101101011111011101101111001101101011111101111;
                    10: level_vec_out = 100'b1111111001111101101011001010111101101011100111100101010101101011111011101101111001101101011111101111;
                    11: level_vec_out = 100'b1111111001111101101011001010111101101011100111100101010101101011111011101111111001101101011111101111;
                    12: level_vec_out = 100'b1111111001111101101011001010111101101011100111100101010101101011111011101111111001101101011111101111;
                    13: level_vec_out = 100'b1111111001111101101011001010111101111011100111100101010101101011111011101111111001101111011111101111;
                    14: level_vec_out = 100'b1111111001111101101011001010111101111011100111110101010101101011111011101111111001101111111111101111;
                    15: level_vec_out = 100'b1111111001111101111011001010111101111011100111110101010111101111111011101111111001111111111111101111;
                    16: level_vec_out = 100'b1111111011111101111011111010111101111111100111110101010111101111111011101111111011111111111111111111;
                    17: level_vec_out = 100'b1111111011111111111011111010111101111111110111110101010111101111111011101111111011111111111111111111;
                    18: level_vec_out = 100'b1111111011111111111011111010111101111111110111110101010111101111111011111111111111111111111111111111;
                    19: level_vec_out = 100'b1111111011111111111011111010111101111111110111110101010111101111111011111111111111111111111111111111;
                    20: level_vec_out = 100'b1111111011111111111011111011111101111111111111110101010111101111111011111111111111111111111111111111;
                    21: level_vec_out = 100'b1111111011111111111011111011111101111111111111110101010111101111111011111111111111111111111111111111;
                    22: level_vec_out = 100'b1111111011111111111011111011111101111111111111110101010111101111111011111111111111111111111111111111;
                    23: level_vec_out = 100'b1111111011111111111011111011111101111111111111110101110111101111111011111111111111111111111111111111;
                    24: level_vec_out = 100'b1111111011111111111011111111111101111111111111110101110111101111111011111111111111111111111111111111;
                    25: level_vec_out = 100'b1111111011111111111011111111111101111111111111110101111111111111111011111111111111111111111111111111;
                    26: level_vec_out = 100'b1111111011111111111011111111111101111111111111110111111111111111111011111111111111111111111111111111;
                    27: level_vec_out = 100'b1111111111111111111111111111111101111111111111110111111111111111111011111111111111111111111111111111;
                    28: level_vec_out = 100'b1111111111111111111111111111111111111111111111110111111111111111111011111111111111111111111111111111;
                    29: level_vec_out = 100'b1111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111;
                endcase
            end
            4: begin
                case (frame_id)
                    0: level_vec_out = 100'b0100000110110111001011000001101001001101110001001101011111001110000011011111000110110001011010011111;
                    1: level_vec_out = 100'b0100000110110111001011000001101001001101110001001101011111001110000011011111000110110001011111011111;
                    2: level_vec_out = 100'b0100000110110111001011000001101101001101110001001101011111001110000011011111000110110001011111011111;
                    3: level_vec_out = 100'b0100000110110111101011000001101101001101110001001101011111001110000011011111000110110001011111011111;
                    4: level_vec_out = 100'b0100000110110111101011000101101101001101110001001101011111001110000011011111000110110001011111011111;
                    5: level_vec_out = 100'b0100000110110111101011000101101101001101110001001101011111001110000011011111000110110001011111011111;
                    6: level_vec_out = 100'b0100000110110111101011000101101101001101110001001101011111101110000011011111001110110001011111011111;
                    7: level_vec_out = 100'b0100010110110111101011000101101101001101110001001111011111101110000011011111001110110001011111011111;
                    8: level_vec_out = 100'b1100010110110111101011000101101101001101110001001111111111101110100011011111001110110001011111111111;
                    9: level_vec_out = 100'b1100010110110111101011000101101101001101110001001111111111101110100011011111001110110001011111111111;
                    10: level_vec_out = 100'b1100010110110111101011000101101101001101110001001111111111101110101011011111001110110001011111111111;
                    11: level_vec_out = 100'b1100010110110111101011000101101101001101110001001111111111101110101011011111001110110001011111111111;
                    12: level_vec_out = 100'b1100010110110111101011000101101101001101110001001111111111101110101011011111101110110001011111111111;
                    13: level_vec_out = 100'b1100010110110111101011000101101101001101110001001111111111101110101011011111101110110001011111111111;
                    14: level_vec_out = 100'b1100110110110111101011000101101101011101110001001111111111101110101011011111101110110101011111111111;
                    15: level_vec_out = 100'b1100110110110111101011000101101101011101110001101111111111101110101011011111101110110101011111111111;
                    16: level_vec_out = 100'b1101110110110111101011000101101101011101110001101111111111101110101011011111101110110101011111111111;
                    17: level_vec_out = 100'b1101110110110111101111000101101101011101110001101111111111101111101011011111101111110101011111111111;
                    18: level_vec_out = 100'b1101110110110111101111000101101101011101110001101111111111101111101011011111101111110101011111111111;
                    19: level_vec_out = 100'b1101110110111111101111000101101101011101110001101111111111101111101011011111101111110101011111111111;
                    20: level_vec_out = 100'b1111110110111111101111000101101101011101111001101111111111101111111011011111101111110101011111111111;
                    21: level_vec_out = 100'b1111110110111111101111100101111101011101111101101111111111101111111011011111101111111101011111111111;
                    22: level_vec_out = 100'b1111111110111111101111100101111101011101111101101111111111111111111011011111101111111101111111111111;
                    23: level_vec_out = 100'b1111111110111111101111110101111101011101111101111111111111111111111011011111101111111101111111111111;
                    24: level_vec_out = 100'b1111111110111111101111110111111101011111111101111111111111111111111011011111101111111101111111111111;
                    25: level_vec_out = 100'b1111111110111111101111110111111101011111111101111111111111111111111011011111101111111111111111111111;
                    26: level_vec_out = 100'b1111111110111111111111110111111101011111111101111111111111111111111011011111111111111111111111111111;
                    27: level_vec_out = 100'b1111111110111111111111110111111101111111111101111111111111111111111011011111111111111111111111111111;
                    28: level_vec_out = 100'b1111111110111111111111110111111101111111111101111111111111111111111011011111111111111111111111111111;
                    29: level_vec_out = 100'b1111111110111111111111110111111101111111111101111111111111111111111011011111111111111111111111111111;
                endcase
            end
            5: begin
                case (frame_id)
                    0: level_vec_out = 100'b1010110000010000110100010000101110010100010010000000001110011100001101011010000000000000010000001000;
                    1: level_vec_out = 100'b1010110000010000110100010000101110010100010010000000001110011101001101011010000000000100010001001000;
                    2: level_vec_out = 100'b1010110000010000111100110000101110010100010010000000011110011101001111011010000000100100010001001000;
                    3: level_vec_out = 100'b1010110000010000111100110000101110010100010010000000011110011101001111011010000000100100010001001000;
                    4: level_vec_out = 100'b1010110000010000111100110000101110010110010010000000011110011101001111011010100000100100010001001000;
                    5: level_vec_out = 100'b1010110000010000111100110000101110010110010010000000111110011101001111011010100000100101010011001000;
                    6: level_vec_out = 100'b1010110000010000111100110001101110010110010010010000111110011101001111011010100000100101010011001000;
                    7: level_vec_out = 100'b1010110000010000111100110001101110010110010110110000111110011101001111011010100000100101010011001100;
                    8: level_vec_out = 100'b1010110000010000111100110001101110010110010111110000111110011101001111011010110100100101010011001101;
                    9: level_vec_out = 100'b1010110001110000111101110001101110010110010111110000111110011101001111011010110101100101110011001101;
                    10: level_vec_out = 100'b1010110101110001111111110001101110010110010111110000111110011101001111011010110101100101110011001101;
                    11: level_vec_out = 100'b1010110111110001111111110001101110010110010111110000111111011101101111011010110101110101110011001101;
                    12: level_vec_out = 100'b1010110111110001111111110001101110010110010111110000111111011101101111011010110101110101110111001101;
                    13: level_vec_out = 100'b1010110111110001111111110001101110010110010111110000111111011101101111011010111101110111110111001101;
                    14: level_vec_out = 100'b1010110111110101111111110001101110110110010111110000111111011101101111011010111101110111110111001101;
                    15: level_vec_out = 100'b1010110111110101111111110001101110110110011111110000111111011101101111011010111101110111110111001101;
                    16: level_vec_out = 100'b1010110111110101111111110001101110110110011111110000111111011101101111011010111101110111110111001101;
                    17: level_vec_out = 100'b1010110111110101111111110001101110110111011111110000111111011101101111011010111101110111110111001101;
                    18: level_vec_out = 100'b1010110111111101111111111001101110110111011111110000111111011101101111011010111101110111110111001101;
                    19: level_vec_out = 100'b1010110111111111111111111001101110110111011111110000111111011101101111011110111101110111110111001101;
                    20: level_vec_out = 100'b1010110111111111111111111001101110110111011111110001111111011101101111011111111101110111110111001101;
                    21: level_vec_out = 100'b1011110111111111111111111001101110110111011111110001111111011101101111011111111101110111110111101101;
                    22: level_vec_out = 100'b1111110111111111111111111101101110110111011111110001111111011101101111111111111101110111110111101111;
                    23: level_vec_out = 100'b1111110111111111111111111101101110110111011111110001111111011101101111111111111101110111110111101111;
                    24: level_vec_out = 100'b1111110111111111111111111101101110110111011111110001111111111101101111111111111111111111110111101111;
                    25: level_vec_out = 100'b1111110111111111111111111101111110110111011111110001111111111101101111111111111111111111110111101111;
                    26: level_vec_out = 100'b1111110111111111111111111111111110110111011111110001111111111101101111111111111111111111110111101111;
                    27: level_vec_out = 100'b1111110111111111111111111111111110110111011111110001111111111101101111111111111111111111110111101111;
                    28: level_vec_out = 100'b1111110111111111111111111111111111111111111111110001111111111101101111111111111111111111110111101111;
                    29: level_vec_out = 100'b1111110111111111111111111111111111111111111111110101111111111101101111111111111111111111111111101111;
                endcase
            end
            6: begin
                case (frame_id)
                    0: level_vec_out = 100'b1110101011000011110010111111010110110111111111111101000101111100100100100011010011101111111000011111;
                    1: level_vec_out = 100'b1110111011000011110010111111010110110111111111111101000101111100100100100011010011101111111000011111;
                    2: level_vec_out = 100'b1110111011000111110010111111010110110111111111111101000101111100100100100011010011101111111000011111;
                    3: level_vec_out = 100'b1110111011100111110010111111010110110111111111111101010101111100100100100011010011101111111000011111;
                    4: level_vec_out = 100'b1110111011100111110010111111010110110111111111111101010101111100100100100011010011101111111000011111;
                    5: level_vec_out = 100'b1110111011100111110010111111010110110111111111111101010101111100100101100011011011101111111000011111;
                    6: level_vec_out = 100'b1110111011101111110010111111010110110111111111111101010101111100100101101011011011101111111000011111;
                    7: level_vec_out = 100'b1110111011101111110110111111010110110111111111111101010101111101100101101011011011101111111000011111;
                    8: level_vec_out = 100'b1110111011101111110110111111010110110111111111111101010101111101101101101011011011101111111000011111;
                    9: level_vec_out = 100'b1110111011101111110110111111010110110111111111111101010101111101101101101011011011111111111000011111;
                    10: level_vec_out = 100'b1110111011101111110110111111010110110111111111111101010101111101101101101011011011111111111001011111;
                    11: level_vec_out = 100'b1110111011101111110110111111010110110111111111111101010101111101101101111011011011111111111001011111;
                    12: level_vec_out = 100'b1110111011101111110110111111010110110111111111111101010101111111101101111011011011111111111001011111;
                    13: level_vec_out = 100'b1110111111111111110110111111010110110111111111111101010101111111101101111011011011111111111001011111;
                    14: level_vec_out = 100'b1110111111111111110110111111010110110111111111111101010101111111101111111011011011111111111001011111;
                    15: level_vec_out = 100'b1110111111111111110110111111010110110111111111111101010101111111101111111011011011111111111001111111;
                    16: level_vec_out = 100'b1110111111111111110110111111010110110111111111111101010101111111101111111011011011111111111001111111;
                    17: level_vec_out = 100'b1110111111111111110110111111010110110111111111111101010101111111101111111011011011111111111001111111;
                    18: level_vec_out = 100'b1110111111111111110110111111010110110111111111111101110101111111101111111011011011111111111001111111;
                    19: level_vec_out = 100'b1110111111111111110110111111010110110111111111111101110101111111101111111011011011111111111001111111;
                    20: level_vec_out = 100'b1110111111111111110110111111010110110111111111111101110101111111101111111011011011111111111001111111;
                    21: level_vec_out = 100'b1110111111111111110110111111010110110111111111111101110101111111101111111011011011111111111011111111;
                    22: level_vec_out = 100'b1110111111111111110111111111010110110111111111111101110101111111111111111111011111111111111011111111;
                    23: level_vec_out = 100'b1110111111111111110111111111010110110111111111111101110111111111111111111111011111111111111011111111;
                    24: level_vec_out = 100'b1110111111111111111111111111010110110111111111111101110111111111111111111111011111111111111011111111;
                    25: level_vec_out = 100'b1110111111111111111111111111010110111111111111111101110111111111111111111111011111111111111011111111;
                    26: level_vec_out = 100'b1110111111111111111111111111010110111111111111111101110111111111111111111111011111111111111111111111;
                    27: level_vec_out = 100'b1110111111111111111111111111010110111111111111111101111111111111111111111111011111111111111111111111;
                    28: level_vec_out = 100'b1111111111111111111111111111010110111111111111111111111111111111111111111111111111111111111111111111;
                    29: level_vec_out = 100'b1111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111;
                endcase
            end
            7: begin
                case (frame_id)
                    0: level_vec_out = 100'b0001111000101111110100011111100001000110011000010101100111100101100111010101011001011100001001111101;
                    1: level_vec_out = 100'b0101111000101111110100011111100001000110011000010101100111100101100111010101011001011100001001111111;
                    2: level_vec_out = 100'b0101111000101111110100011111100111000110011000010101100111100101100111010101011001011100001001111111;
                    3: level_vec_out = 100'b0101111000101111110100011111100111000110011000010101100111100101100111010101111001011100001001111111;
                    4: level_vec_out = 100'b0101111000101111110100011111100111000110011000010101100111100101100111010101111001011100001001111111;
                    5: level_vec_out = 100'b0111111000101111110100011111100111000110011000010101100111100101110111010101111001011100001001111111;
                    6: level_vec_out = 100'b0111111000101111110100011111100111000110011000010101100111100101110111010101111001011100001001111111;
                    7: level_vec_out = 100'b0111111000101111110100011111100111100110011000010101100111100101110111010101111101011100001001111111;
                    8: level_vec_out = 100'b0111111001101111110100011111100111100110011000010101100111100101110111010101111101011100001001111111;
                    9: level_vec_out = 100'b0111111001101111110100011111100111110110011000010101100111100101110111010101111101011100001001111111;
                    10: level_vec_out = 100'b0111111001101111110100011111100111110110011000010101100111100101110111010101111101011100101001111111;
                    11: level_vec_out = 100'b0111111001101111110100011111100111111110011010110101100111110101110111010101111101011100101001111111;
                    12: level_vec_out = 100'b0111111001101111110100011111100111111110011010111101100111110101110111010101111101011100101001111111;
                    13: level_vec_out = 100'b0111111001101111110100011111100111111110011010111101100111111101110111010101111101011101101001111111;
                    14: level_vec_out = 100'b0111111001101111110100011111100111111110011010111101100111111101110111010101111101011101101011111111;
                    15: level_vec_out = 100'b0111111001101111110100011111100111111110011010111101100111111101111111010101111101011101101011111111;
                    16: level_vec_out = 100'b0111111001101111110100011111100111111110011011111101100111111101111111110101111101011101101011111111;
                    17: level_vec_out = 100'b0111111001101111110100111111100111111110011011111101100111111101111111111101111101011101101011111111;
                    18: level_vec_out = 100'b0111111001101111110100111111100111111110011011111101100111111101111111111101111101011101101011111111;
                    19: level_vec_out = 100'b0111111001101111110101111111100111111110011011111101100111111101111111111111111101011101101011111111;
                    20: level_vec_out = 100'b0111111001101111110111111111100111111110011011111101100111111101111111111111111101011101101011111111;
                    21: level_vec_out = 100'b1111111001101111110111111111100111111110011011111101100111111101111111111111111101011101101011111111;
                    22: level_vec_out = 100'b1111111001101111110111111111100111111110011011111101100111111101111111111111111101011101101011111111;
                    23: level_vec_out = 100'b1111111001101111110111111111100111111110111011111101100111111101111111111111111101011101101011111111;
                    24: level_vec_out = 100'b1111111001101111110111111111100111111111111111111101100111111101111111111111111101011101101011111111;
                    25: level_vec_out = 100'b1111111001111111110111111111100111111111111111111101100111111101111111111111111101011111101011111111;
                    26: level_vec_out = 100'b1111111101111111110111111111100111111111111111111101100111111101111111111111111101111111101011111111;
                    27: level_vec_out = 100'b1111111101111111110111111111101111111111111111111101101111111101111111111111111101111111101011111111;
                    28: level_vec_out = 100'b1111111101111111111111111111111111111111111111111111111111111101111111111111111101111111111011111111;
                    29: level_vec_out = 100'b1111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111011111111;
                endcase
            end
            8: begin
                case (frame_id)
                    0: level_vec_out = 100'b0011110000111111001000001111100011100011110010110101000010001111110010000110100001101011100001010000;
                    1: level_vec_out = 100'b0011110000111111001000011111100011100011110010110101000010001111110010000110100001101011100001010000;
                    2: level_vec_out = 100'b0011110000111111001000011111100011100011110010110101000010001111110010000110100001101011100001010000;
                    3: level_vec_out = 100'b0011110000111111001000011111101111100011110010110101001010001111110010000110100001101011100001010000;
                    4: level_vec_out = 100'b1011110000111111001000011111101111100011110010110101001010001111110010000110100001101011100001010101;
                    5: level_vec_out = 100'b1011110000111111001000011111101111100011110010110101001010001111110010000110100001101011100001010101;
                    6: level_vec_out = 100'b1011110000111111001000011111101111100011111010110101001010001111110010000110100001101011100001010101;
                    7: level_vec_out = 100'b1011110000111111001000011111101111100011111010111101001010001111110010000110100001101011100001010101;
                    8: level_vec_out = 100'b1011110000111111001000011111101111100011111010111101001010001111110010000110100001101011101101010101;
                    9: level_vec_out = 100'b1011110000111111001100011111101111100011111010111101001010011111110110000110100001101011101101010101;
                    10: level_vec_out = 100'b1011110001111111001100011111101111100011111011111101001110011111110110000110111001101011101101110101;
                    11: level_vec_out = 100'b1011110001111111001100011111101111100011111011111101001110011111110110000110111001101011101101110101;
                    12: level_vec_out = 100'b1011110001111111001100011111101111100011111011111101001110011111110110001110111001111011111101110101;
                    13: level_vec_out = 100'b1011110001111111001100011111101111100011111011111101001110011111110111001110111001111011111111110101;
                    14: level_vec_out = 100'b1011110001111111001100011111101111100011111011111101001110011111110111001110111001111011111111110101;
                    15: level_vec_out = 100'b1011110001111111001101011111101111110011111111111101011110011111110111011110111001111011111111110101;
                    16: level_vec_out = 100'b1111110011111111001101011111101111110011111111111101011110011111110111011110111101111011111111110101;
                    17: level_vec_out = 100'b1111110111111111001101111111101111110011111111111101011110011111110111011110111101111011111111110101;
                    18: level_vec_out = 100'b1111110111111111001101111111101111110011111111111101011110011111110111011110111101111011111111110101;
                    19: level_vec_out = 100'b1111110111111111001101111111101111110011111111111101011110011111110111011110111101111011111111110101;
                    20: level_vec_out = 100'b1111110111111111001101111111111111110011111111111101011110111111110111011110111101111011111111110101;
                    21: level_vec_out = 100'b1111110111111111001101111111111111110011111111111101111111111111111111011111111101111011111111110101;
                    22: level_vec_out = 100'b1111110111111111001101111111111111111011111111111101111111111111111111011111111101111011111111110101;
                    23: level_vec_out = 100'b1111110111111111001101111111111111111011111111111111111111111111111111011111111111111111111111110101;
                    24: level_vec_out = 100'b1111110111111111001101111111111111111011111111111111111111111111111111011111111111111111111111110101;
                    25: level_vec_out = 100'b1111110111111111001101111111111111111011111111111111111111111111111111011111111111111111111111110101;
                    26: level_vec_out = 100'b1111110111111111101101111111111111111111111111111111111111111111111111011111111111111111111111110101;
                    27: level_vec_out = 100'b1111111111111111101101111111111111111111111111111111111111111111111111011111111111111111111111110101;
                    28: level_vec_out = 100'b1111111111111111101101111111111111111111111111111111111111111111111111011111111111111111111111110101;
                    29: level_vec_out = 100'b1111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111110101;
                endcase
            end
            9: begin
                case (frame_id)
                    0: level_vec_out = 100'b1001101110101110010110101110101101010101010011011111011000110100011001010100010000110010001101101010;
                    1: level_vec_out = 100'b1001101110101110010110101110101101010101010011011111111000110110011001010100010000110010001101101010;
                    2: level_vec_out = 100'b1001101110101110010110101110101101010101010011011111111000110110011001010100011000110011001101101010;
                    3: level_vec_out = 100'b1101111110101110010110101110101101010101010011011111111000110111011001110100011000110011001101101010;
                    4: level_vec_out = 100'b1101111110101110010111101110101101010101010011011111111000110111011001110100011010110011001101101010;
                    5: level_vec_out = 100'b1101111110101110110111101110101101010101010011011111111000110111011001110100011010110011001101111010;
                    6: level_vec_out = 100'b1101111110101110110111101110101101010101010011011111111100110111011001110100011010110011001101111010;
                    7: level_vec_out = 100'b1101111110101110110111101110101101010101010011011111111110110111011001110100011010110011001101111010;
                    8: level_vec_out = 100'b1101111110101110110111101110101101010101010011011111111110110111011001110100011110110011001101111010;
                    9: level_vec_out = 100'b1101111110101110110111101110101101010101010011011111111110110111011011110100011110110011001101111010;
                    10: level_vec_out = 100'b1101111110101110110111101110101101010101010011011111111110110111011011110100011110110011001101111010;
                    11: level_vec_out = 100'b1101111110101110110111101110101101010101010011011111111110110111011011110100011110110011001101111110;
                    12: level_vec_out = 100'b1101111110101110110111101110101101010101010111011111111110110111011111110100011110110011001101111110;
                    13: level_vec_out = 100'b1101111110101110110111111110101101010101010111111111111110110111011111110110011110110011001101111110;
                    14: level_vec_out = 100'b1101111110101110110111111110101101010101010111111111111110110111011111110110011111110011011101111110;
                    15: level_vec_out = 100'b1101111110101110110111111110111101010101010111111111111110110111011111110110011111110011011101111110;
                    16: level_vec_out = 100'b1101111110101110110111111110111101010101010111111111111110110111011111110110011111110011011101111110;
                    17: level_vec_out = 100'b1101111110101110110111111110111111011101010111111111111110110111011111110110011111110011011101111110;
                    18: level_vec_out = 100'b1101111111101110110111111110111111011101010111111111111110110111011111110110011111110111111101111110;
                    19: level_vec_out = 100'b1101111111101110110111111110111111011101010111111111111110110111111111110110011111111111111101111110;
                    20: level_vec_out = 100'b1101111111101110110111111110111111011101010111111111111110110111111111110110011111111111111101111110;
                    21: level_vec_out = 100'b1111111111101110110111111110111111011101010111111111111110110111111111110111011111111111111101111110;
                    22: level_vec_out = 100'b1111111111101110110111111110111111111101010111111111111110110111111111110111011111111111111101111110;
                    23: level_vec_out = 100'b1111111111101110110111111110111111111101010111111111111110110111111111110111011111111111111101111110;
                    24: level_vec_out = 100'b1111111111101110110111111110111111111101010111111111111110110111111111110111011111111111111111111111;
                    25: level_vec_out = 100'b1111111111111110110111111110111111111101010111111111111110110111111111110111011111111111111111111111;
                    26: level_vec_out = 100'b1111111111111110110111111110111111111111010111111111111110110111111111110111011111111111111111111111;
                    27: level_vec_out = 100'b1111111111111110110111111111111111111111110111111111111111110111111111110111011111111111111111111111;
                    28: level_vec_out = 100'b1111111111111110110111111111111111111111110111111111111111110111111111110111011111111111111111111111;
                    29: level_vec_out = 100'b1111111111111110110111111111111111111111110111111111111111110111111111110111011111111111111111111111;
                endcase
            end
        endcase
    end
endmodule