----
 -- @file level_hvec_gen_hdl.hpp
 -- @brief This script generates HDL code for generating high-dimensional LEVEL vectors.
 -- It is a novel method; for more information, please refer to our paper.
 --
 -- @author Saeid Jamili and Marco Angioli
 -- @note Author names are listed in alphabetical order.
 -- @email <saeid.jamili@uniroma1.it>
 -- @email <marco.angioli@uniroma1.it>
 --
 -- @contributors
 --
 -- @date Created: 24th July 2023
 -- @date Last Updated: 23th August 2023
 --
 -- @version 1.0.0
 --
 -- @institute Sapienza University of Rome
 -- @cite https://doi.org/10.xxxx/yyyyy
 --
 -- @section DEPENDENCIES
 -- - Dependency1: Description or version details.
 -- - Dependency2: Description or version details.
 --
 -- @section LICENSE
 -- This file is part of the Aeneas HyperCompute Platform.
 --
 -- Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 --
 -- @section CHANGELOG
 -- @version 1.0.0-dev - 23th August 2023
 -- - Initial release
 --
 -- @todo
 -- - Complete level vector generator function
 -- - Add training
 --
 -- @see
 -- -
 -- -
 -- -
 --
 --

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity level_vec_gen is
    Port ( level_vec_out : out  STD_LOGIC_VECTOR (63 downto 0);
           frame_index : in  STD_LOGIC_VECTOR (2 downto 0);
           frame_id : in  STD_LOGIC_VECTOR (4 downto 0));
end level_vec_gen;

architecture Behavioral of level_vec_gen is
begin
    process (frame_index, frame_id)
    begin
        -- Update this function to match your requirements
        case frame_index is
            when "000" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1010101110011010000001100011010101000001111011110100100001001001";
                    when "00001" => level_vec_out <= "1010101110111010000001100011010101000001111011110100100001001001";
                    when "00010" => level_vec_out <= "1010101110111010000001100111011101000001111011110100100001001001";
                    when "00011" => level_vec_out <= "1010101110111010000001100111011101000001111011110100100011001001";
                    when "00100" => level_vec_out <= "1010101110111010000001100111011101000001111011110100100011001001";
                    when "00101" => level_vec_out <= "1010101110111010000001100111011101000001111011110100100011001001";
                    when "00110" => level_vec_out <= "1010101110111010000001100111011101000001111011110100110011001001";
                    when "00111" => level_vec_out <= "1010101110111010000001100111011101000001111011110100110011001001";
                    when "01000" => level_vec_out <= "1010101110111010100001101111011101000001111011110101110011001001";
                    when "01001" => level_vec_out <= "1010101110111010100001101111011101000001111011110101110011001001";
                    when "01010" => level_vec_out <= "1110101110111010100001101111011101000001111011110101110011001001";
                    when "01011" => level_vec_out <= "1110101110111010100001101111011101001001111011110101110011001001";
                    when "01100" => level_vec_out <= "1110101110111010100001101111011101001011111011110101110011001001";
                    when "01101" => level_vec_out <= "1110101110111010100001101111011101001011111011110101110011001001";
                    when "01110" => level_vec_out <= "1110101110111010110001101111111101001011111011110101111011001001";
                    when "01111" => level_vec_out <= "1110101110111010110011101111111101001011111011110101111011001001";
                    when "10000" => level_vec_out <= "1110101110111010110011111111111101001011111011110101111011001001";
                    when "10001" => level_vec_out <= "1110101110111010110011111111111101001111111011110101111011001001";
                    when "10010" => level_vec_out <= "1111101110111010110011111111111101001111111011110101111011001001";
                    when "10011" => level_vec_out <= "1111101110111010110011111111111101001111111011110101111011101001";
                    when "10100" => level_vec_out <= "1111101110111110110011111111111101001111111011110101111011111001";
                    when "10101" => level_vec_out <= "1111101110111110110011111111111101001111111111110101111011111001";
                    when "10110" => level_vec_out <= "1111101110111110110011111111111101001111111111110101111011111001";
                    when "10111" => level_vec_out <= "1111101110111111110011111111111101001111111111110111111011111001";
                    when "11000" => level_vec_out <= "1111101110111111110011111111111101001111111111110111111011111001";
                    when "11001" => level_vec_out <= "1111101111111111110011111111111101001111111111110111111011111001";
                    when "11010" => level_vec_out <= "1111101111111111110011111111111101001111111111110111111011111001";
                    when "11011" => level_vec_out <= "1111101111111111111111111111111101101111111111110111111011111001";
                    when "11100" => level_vec_out <= "1111101111111111111111111111111101101111111111111111111011111101";
                    when "11101" => level_vec_out <= "1111101111111111111111111111111111101111111111111111111011111101";
                    when "11110" => level_vec_out <= "1111101111111111111111111111111111101111111111111111111011111101";
                    when "11111" => level_vec_out <= "1111101111111111111111111111111111111111111111111111111011111111";
                when others => null;
                end case;
            when "001" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0101000101111001100010111000001111001010001110010010111001001110";
                    when "00001" => level_vec_out <= "0101000101111001100010111000001111001010011110010010111001001110";
                    when "00010" => level_vec_out <= "0101000101111001100010111000001111001010011110010010111001001110";
                    when "00011" => level_vec_out <= "0101000101111001100010111010001111001010011111010010111001001110";
                    when "00100" => level_vec_out <= "0101000101111001100010111010001111001010011111010010111001001110";
                    when "00101" => level_vec_out <= "0101100101111001110010111010001111001010011111010010111001001110";
                    when "00110" => level_vec_out <= "0101100101111001110010111010001111001010011111110010111001001110";
                    when "00111" => level_vec_out <= "0101100101111001110010111010001111001010011111110010111001101111";
                    when "01000" => level_vec_out <= "0101100101111001110010111010001111001010011111110010111001101111";
                    when "01001" => level_vec_out <= "0101100101111001110110111010001111101010011111110010111001111111";
                    when "01010" => level_vec_out <= "0101100101111001110110111010001111101010011111110010111001111111";
                    when "01011" => level_vec_out <= "0101100101111001110110111010001111101010011111110010111001111111";
                    when "01100" => level_vec_out <= "0111100101111001110110111010001111101010011111110110111001111111";
                    when "01101" => level_vec_out <= "0111100101111001110110111010001111101011011111110110111101111111";
                    when "01110" => level_vec_out <= "0111100101111001110110111010001111101011011111110110111101111111";
                    when "01111" => level_vec_out <= "0111100101111001110110111010001111101011011111110110111101111111";
                    when "10000" => level_vec_out <= "0111110101111001110110111010011111101011011111110110111101111111";
                    when "10001" => level_vec_out <= "0111110101111001110110111010111111101011011111110110111101111111";
                    when "10010" => level_vec_out <= "0111110101111001110111111010111111101011011111110110111101111111";
                    when "10011" => level_vec_out <= "0111110101111001110111111010111111101011011111110110111101111111";
                    when "10100" => level_vec_out <= "0111110101111001110111111010111111101011011111110110111101111111";
                    when "10101" => level_vec_out <= "0111110101111011110111111010111111101011011111110110111101111111";
                    when "10110" => level_vec_out <= "0111111101111011111111111010111111101011011111110110111101111111";
                    when "10111" => level_vec_out <= "0111111101111111111111111010111111101011011111110110111111111111";
                    when "11000" => level_vec_out <= "1111111101111111111111111010111111101011011111110110111111111111";
                    when "11001" => level_vec_out <= "1111111101111111111111111010111111101011011111110110111111111111";
                    when "11010" => level_vec_out <= "1111111101111111111111111010111111111011011111110111111111111111";
                    when "11011" => level_vec_out <= "1111111111111111111111111010111111111111011111110111111111111111";
                    when "11100" => level_vec_out <= "1111111111111111111111111110111111111111011111110111111111111111";
                    when "11101" => level_vec_out <= "1111111111111111111111111110111111111111111111110111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "010" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1100110010010110001110110001110111010100111110101000100100010001";
                    when "00001" => level_vec_out <= "1100110010010110001110110001110111010100111110101000100100010001";
                    when "00010" => level_vec_out <= "1100110110010110001110110001110111010100111110101000100100010001";
                    when "00011" => level_vec_out <= "1100110110010110001110110001110111010100111110111010100100010001";
                    when "00100" => level_vec_out <= "1100110110010110001110110001110111010100111110111010100100010001";
                    when "00101" => level_vec_out <= "1100110110010110001110110011110111010110111110111010100100010001";
                    when "00110" => level_vec_out <= "1100110110010110001110110011110111110110111110111010101100010001";
                    when "00111" => level_vec_out <= "1101110110010110001110111011110111110110111110111010101100010001";
                    when "01000" => level_vec_out <= "1101110110010110001110111011110111110110111110111010101100010001";
                    when "01001" => level_vec_out <= "1101110110010110001110111011110111110110111110111010101100010001";
                    when "01010" => level_vec_out <= "1101110110010110001110111111110111110110111110111010101101010011";
                    when "01011" => level_vec_out <= "1111110110010110101110111111110111110110111110111110101101010011";
                    when "01100" => level_vec_out <= "1111110110010110101110111111110111110110111110111110101101010011";
                    when "01101" => level_vec_out <= "1111110110011110101110111111110111110110111110111110101101010011";
                    when "01110" => level_vec_out <= "1111110110011110101110111111110111110110111110111111101101110011";
                    when "01111" => level_vec_out <= "1111110110011110101110111111110111110110111110111111101101110011";
                    when "10000" => level_vec_out <= "1111110110011110101110111111110111110110111110111111101101110011";
                    when "10001" => level_vec_out <= "1111110110111110101110111111110111110110111110111111101101110011";
                    when "10010" => level_vec_out <= "1111110110111110101110111111110111110110111110111111101101111011";
                    when "10011" => level_vec_out <= "1111110110111110101110111111111111110111111110111111101111111011";
                    when "10100" => level_vec_out <= "1111110110111111111110111111111111110111111110111111101111111011";
                    when "10101" => level_vec_out <= "1111110110111111111110111111111111110111111110111111101111111011";
                    when "10110" => level_vec_out <= "1111110110111111111110111111111111110111111111111111111111111011";
                    when "10111" => level_vec_out <= "1111111110111111111111111111111111111111111111111111111111111011";
                    when "11000" => level_vec_out <= "1111111110111111111111111111111111111111111111111111111111111011";
                    when "11001" => level_vec_out <= "1111111110111111111111111111111111111111111111111111111111111011";
                    when "11010" => level_vec_out <= "1111111110111111111111111111111111111111111111111111111111111011";
                    when "11011" => level_vec_out <= "1111111110111111111111111111111111111111111111111111111111111011";
                    when "11100" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111011";
                    when "11101" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111011";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111011";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111011";
                when others => null;
                end case;
            when "011" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1101010011000100101111110011110110101101001001010001010010001100";
                    when "00001" => level_vec_out <= "1101010011000100101111110011110110101101101001010001010010001100";
                    when "00010" => level_vec_out <= "1101010011000100101111111011110110101101101001010001010010001100";
                    when "00011" => level_vec_out <= "1101010011000100101111111011110110101101101001010001010010001100";
                    when "00100" => level_vec_out <= "1101010011000100101111111011110110101101101001010001010010001101";
                    when "00101" => level_vec_out <= "1111010011000100101111111011110110101101101001010001010010001101";
                    when "00110" => level_vec_out <= "1111010011000100101111111011110110101101101001010001010010001101";
                    when "00111" => level_vec_out <= "1111010011010100101111111011110110101101101001010001010010001101";
                    when "01000" => level_vec_out <= "1111010011010100101111111011110110111101101001010001010010001101";
                    when "01001" => level_vec_out <= "1111010111010100101111111011110110111101101011010001010010001101";
                    when "01010" => level_vec_out <= "1111010111010100101111111011111110111101101011010001010010011101";
                    when "01011" => level_vec_out <= "1111010111010100101111111011111111111101101011010001010010011101";
                    when "01100" => level_vec_out <= "1111010111010100101111111011111111111101101011010001010110011101";
                    when "01101" => level_vec_out <= "1111010111010100101111111011111111111101101011010001010110011101";
                    when "01110" => level_vec_out <= "1111010111110110101111111011111111111101101011010001010110011101";
                    when "01111" => level_vec_out <= "1111010111110110101111111011111111111101101011010001010110011101";
                    when "10000" => level_vec_out <= "1111010111110110101111111011111111111101101011110001010110011101";
                    when "10001" => level_vec_out <= "1111010111110110101111111011111111111101101011110001010110011101";
                    when "10010" => level_vec_out <= "1111010111110110101111111011111111111111101011110001010110011101";
                    when "10011" => level_vec_out <= "1111010111110110101111111111111111111111101011110001010110011101";
                    when "10100" => level_vec_out <= "1111010111110110101111111111111111111111101011110001010110011101";
                    when "10101" => level_vec_out <= "1111010111110110111111111111111111111111101011110001010110011101";
                    when "10110" => level_vec_out <= "1111010111110111111111111111111111111111101011110101010110011101";
                    when "10111" => level_vec_out <= "1111010111110111111111111111111111111111101011110101010110011101";
                    when "11000" => level_vec_out <= "1111110111110111111111111111111111111111101011110111110110011101";
                    when "11001" => level_vec_out <= "1111110111110111111111111111111111111111101011110111111110011101";
                    when "11010" => level_vec_out <= "1111110111110111111111111111111111111111101111110111111110011101";
                    when "11011" => level_vec_out <= "1111110111110111111111111111111111111111101111110111111110011101";
                    when "11100" => level_vec_out <= "1111110111110111111111111111111111111111111111110111111110111101";
                    when "11101" => level_vec_out <= "1111111111110111111111111111111111111111111111110111111110111101";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111110111101";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111101";
                when others => null;
                end case;
            when "100" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1011100111100001100100010001101110110100000110111010000111111111";
                    when "00001" => level_vec_out <= "1011100111100001100100010001101110110100011110111010000111111111";
                    when "00010" => level_vec_out <= "1011100111110001100100010001101110111100011111111010000111111111";
                    when "00011" => level_vec_out <= "1011100111110001100100010001101110111100011111111010100111111111";
                    when "00100" => level_vec_out <= "1011100111110001100100010001101110111100011111111010100111111111";
                    when "00101" => level_vec_out <= "1011100111110001100100010001101110111100011111111010100111111111";
                    when "00110" => level_vec_out <= "1011100111110001100100010001101110111100011111111010100111111111";
                    when "00111" => level_vec_out <= "1011110111110001100100010001101110111100011111111010100111111111";
                    when "01000" => level_vec_out <= "1011110111110001100100010001101110111100111111111010100111111111";
                    when "01001" => level_vec_out <= "1011110111110001100100110001101110111101111111111010100111111111";
                    when "01010" => level_vec_out <= "1011110111110001100100110011101110111101111111111010100111111111";
                    when "01011" => level_vec_out <= "1011110111110001100100110011111110111101111111111010100111111111";
                    when "01100" => level_vec_out <= "1011110111110101100101110011111110111101111111111010100111111111";
                    when "01101" => level_vec_out <= "1011110111110101100101110011111110111101111111111010100111111111";
                    when "01110" => level_vec_out <= "1011110111110101100101110011111110111101111111111010100111111111";
                    when "01111" => level_vec_out <= "1011110111110101100101110011111110111101111111111010100111111111";
                    when "10000" => level_vec_out <= "1111110111110111100101110011111110111101111111111010100111111111";
                    when "10001" => level_vec_out <= "1111110111110111100101110011111110111101111111111010100111111111";
                    when "10010" => level_vec_out <= "1111110111110111100101110011111111111111111111111010100111111111";
                    when "10011" => level_vec_out <= "1111110111110111100101110011111111111111111111111010100111111111";
                    when "10100" => level_vec_out <= "1111110111110111100101110011111111111111111111111010100111111111";
                    when "10101" => level_vec_out <= "1111110111110111100101110011111111111111111111111110100111111111";
                    when "10110" => level_vec_out <= "1111110111110111100101110011111111111111111111111110101111111111";
                    when "10111" => level_vec_out <= "1111110111110111100101110011111111111111111111111110101111111111";
                    when "11000" => level_vec_out <= "1111110111110111101101110011111111111111111111111110101111111111";
                    when "11001" => level_vec_out <= "1111110111110111101101110011111111111111111111111110111111111111";
                    when "11010" => level_vec_out <= "1111111111111111111101110011111111111111111111111110111111111111";
                    when "11011" => level_vec_out <= "1111111111111111111101110011111111111111111111111110111111111111";
                    when "11100" => level_vec_out <= "1111111111111111111101111011111111111111111111111110111111111111";
                    when "11101" => level_vec_out <= "1111111111111111111111111011111111111111111111111110111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111011111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "101" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0000101001111100010010101011101110011001111100100101001100010110";
                    when "00001" => level_vec_out <= "0000101001111100010010101011101110011001111100100101011100010110";
                    when "00010" => level_vec_out <= "0000101001111100010010101011101110011001111100100101011100010110";
                    when "00011" => level_vec_out <= "0000101001111100010010101011101110011001111100100101011100010110";
                    when "00100" => level_vec_out <= "0000101001111100010011101011101110011001111101100101011100010110";
                    when "00101" => level_vec_out <= "0000101001111100010011101111101110011001111111100101011100010110";
                    when "00110" => level_vec_out <= "0000101001111100010011101111101110011001111111100101011100010110";
                    when "00111" => level_vec_out <= "0000101001111100010011101111101110011001111111100101011100010110";
                    when "01000" => level_vec_out <= "0000101001111100010111101111101110011001111111100101011100010110";
                    when "01001" => level_vec_out <= "0000101001111100010111101111101110011001111111100101011100010110";
                    when "01010" => level_vec_out <= "0000101001111100010111101111101110011001111111100101011100010110";
                    when "01011" => level_vec_out <= "0000101001111100010111101111101110011001111111100101011100010110";
                    when "01100" => level_vec_out <= "0000101001111100010111101111101110011001111111100101011100010110";
                    when "01101" => level_vec_out <= "0001101001111100010111101111101110011001111111100101111100010110";
                    when "01110" => level_vec_out <= "0001101001111100010111101111101110011001111111100101111100010110";
                    when "01111" => level_vec_out <= "0101101001111100010111111111101110011001111111100101111100010110";
                    when "10000" => level_vec_out <= "0111101001111100010111111111101110011001111111100101111100010110";
                    when "10001" => level_vec_out <= "0111111001111100010111111111101110011001111111100111111100010110";
                    when "10010" => level_vec_out <= "0111111001111100011111111111101110111001111111100111111100010110";
                    when "10011" => level_vec_out <= "0111111001111100011111111111101111111001111111100111111100010110";
                    when "10100" => level_vec_out <= "0111111001111110011111111111111111111001111111100111111100010110";
                    when "10101" => level_vec_out <= "0111111011111110011111111111111111111001111111100111111100010110";
                    when "10110" => level_vec_out <= "0111111011111110011111111111111111111001111111100111111100010110";
                    when "10111" => level_vec_out <= "0111111011111110011111111111111111111001111111110111111100010110";
                    when "11000" => level_vec_out <= "0111111011111110011111111111111111111001111111110111111100011111";
                    when "11001" => level_vec_out <= "1111111111111110011111111111111111111101111111110111111100011111";
                    when "11010" => level_vec_out <= "1111111111111110011111111111111111111101111111110111111110011111";
                    when "11011" => level_vec_out <= "1111111111111110011111111111111111111101111111110111111110111111";
                    when "11100" => level_vec_out <= "1111111111111110011111111111111111111101111111110111111110111111";
                    when "11101" => level_vec_out <= "1111111111111110011111111111111111111101111111111111111110111111";
                    when "11110" => level_vec_out <= "1111111111111111011111111111111111111101111111111111111110111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111110111111";
                when others => null;
                end case;
            when "110" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0011000110001011001010010111100001011011110010111110000001011010";
                    when "00001" => level_vec_out <= "0111000110001011001010011111100001011011110010111110000001011010";
                    when "00010" => level_vec_out <= "0111000110001011001010011111100001011011110010111110000001011010";
                    when "00011" => level_vec_out <= "0111000110001011001010011111100001011011110010111110000001011010";
                    when "00100" => level_vec_out <= "0111000110001011001010011111100001011011110010111110000001011011";
                    when "00101" => level_vec_out <= "0111001110001011001010011111100001011011110010111110000001011011";
                    when "00110" => level_vec_out <= "0111101110001011001010111111100001011011110011111110000001011011";
                    when "00111" => level_vec_out <= "0111101110001011001010111111100001011011110011111110000001011111";
                    when "01000" => level_vec_out <= "0111101110001011001010111111100001011011110011111111000001011111";
                    when "01001" => level_vec_out <= "0111101110001011001010111111100001011011110011111111000001011111";
                    when "01010" => level_vec_out <= "0111101110101011001010111111100001011011110011111111000001011111";
                    when "01011" => level_vec_out <= "0111101110101011001010111111100011011111110011111111000001011111";
                    when "01100" => level_vec_out <= "0111101110101011001010111111100011011111110011111111000111011111";
                    when "01101" => level_vec_out <= "0111101110101011001010111111100011011111110011111111100111011111";
                    when "01110" => level_vec_out <= "0111101110101011001010111111100011011111110011111111100111011111";
                    when "01111" => level_vec_out <= "0111101110111011001010111111100011011111111011111111100111011111";
                    when "10000" => level_vec_out <= "0111101110111011001010111111100011011111111111111111100111011111";
                    when "10001" => level_vec_out <= "0111101110111011001010111111100111011111111111111111100111011111";
                    when "10010" => level_vec_out <= "0111101110111011001010111111100111011111111111111111100111011111";
                    when "10011" => level_vec_out <= "0111101110111011001010111111100111111111111111111111100111011111";
                    when "10100" => level_vec_out <= "0111101110111011001010111111100111111111111111111111100111011111";
                    when "10101" => level_vec_out <= "0111101110111011001010111111111111111111111111111111100111011111";
                    when "10110" => level_vec_out <= "0111101110111011001010111111111111111111111111111111100111011111";
                    when "10111" => level_vec_out <= "0111101110111011001010111111111111111111111111111111100111011111";
                    when "11000" => level_vec_out <= "0111101110111011011010111111111111111111111111111111100111011111";
                    when "11001" => level_vec_out <= "0111101110111011011011111111111111111111111111111111100111111111";
                    when "11010" => level_vec_out <= "0111101110111011011011111111111111111111111111111111100111111111";
                    when "11011" => level_vec_out <= "0111101111111011011011111111111111111111111111111111110111111111";
                    when "11100" => level_vec_out <= "0111101111111011011111111111111111111111111111111111110111111111";
                    when "11101" => level_vec_out <= "1111101111111011011111111111111111111111111111111111110111111111";
                    when "11110" => level_vec_out <= "1111101111111111011111111111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111101111111111011111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "111" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0000111011010011101110100100010011100001101100111101111101000110";
                    when "00001" => level_vec_out <= "0000111011010011101110100100010011100001101100111101111101000110";
                    when "00010" => level_vec_out <= "0000111011011011101110100100010011100001101100111101111101000110";
                    when "00011" => level_vec_out <= "0000111011011011101110110100011011100001101100111101111101000110";
                    when "00100" => level_vec_out <= "0001111011011011101110110110011011100001101100111101111111001110";
                    when "00101" => level_vec_out <= "0001111011011011101110110110011011100001101100111101111111001110";
                    when "00110" => level_vec_out <= "0001111011011011101110110110011011100001101100111101111111011110";
                    when "00111" => level_vec_out <= "0001111011011011101110110110011011100001101101111101111111011110";
                    when "01000" => level_vec_out <= "0011111011011011101110110110011011100001101101111101111111011110";
                    when "01001" => level_vec_out <= "0111111011011011101110110110011011100001101101111101111111011110";
                    when "01010" => level_vec_out <= "0111111011011011101110110110011011100001101101111101111111011110";
                    when "01011" => level_vec_out <= "0111111011011011101110110110011011100001101101111101111111011110";
                    when "01100" => level_vec_out <= "0111111011011011101110110110011011100001101101111101111111011110";
                    when "01101" => level_vec_out <= "0111111011011011101110110110011011110001101101111101111111111110";
                    when "01110" => level_vec_out <= "0111111011011011101110110110011011110001111101111101111111111110";
                    when "01111" => level_vec_out <= "1111111011011011101111110111011011110001111101111101111111111110";
                    when "10000" => level_vec_out <= "1111111011011011101111110111011011110001111101111101111111111110";
                    when "10001" => level_vec_out <= "1111111011011011101111110111011011110011111101111101111111111111";
                    when "10010" => level_vec_out <= "1111111011011011101111110111011011110011111101111101111111111111";
                    when "10011" => level_vec_out <= "1111111011011011101111110111111011110011111101111101111111111111";
                    when "10100" => level_vec_out <= "1111111011011011101111110111111011111011111111111101111111111111";
                    when "10101" => level_vec_out <= "1111111011111011101111110111111011111011111111111101111111111111";
                    when "10110" => level_vec_out <= "1111111011111011101111110111111111111011111111111101111111111111";
                    when "10111" => level_vec_out <= "1111111011111011101111110111111111111011111111111101111111111111";
                    when "11000" => level_vec_out <= "1111111011111011101111110111111111111011111111111101111111111111";
                    when "11001" => level_vec_out <= "1111111011111011101111110111111111111011111111111101111111111111";
                    when "11010" => level_vec_out <= "1111111011111111101111110111111111111011111111111101111111111111";
                    when "11011" => level_vec_out <= "1111111011111111101111110111111111111011111111111101111111111111";
                    when "11100" => level_vec_out <= "1111111011111111101111110111111111111011111111111101111111111111";
                    when "11101" => level_vec_out <= "1111111011111111111111110111111111111011111111111111111111111111";
                    when "11110" => level_vec_out <= "1111111011111111111111110111111111111011111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111110111111111111111111111111111111111111111";
                when others => null;
                end case;
            when others => null;
        end case;
    end process;
end Behavioral;