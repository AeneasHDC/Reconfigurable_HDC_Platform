----
 -- @file level_hvec_gen_hdl.hpp
 -- @brief This script generates HDL code for generating high-dimensional LEVEL vectors.
 -- It is a novel method; for more information, please refer to our paper.
 --
 -- @author Saeid Jamili and Marco Angioli
 -- @note Author names are listed in alphabetical order.
 -- @email <saeid.jamili@uniroma1.it>
 -- @email <marco.angioli@uniroma1.it>
 --
 -- @contributors
 --
 -- @date Created: 24th July 2023
 -- @date Last Updated: 23th August 2023
 --
 -- @version 1.0.0
 --
 -- @institute Sapienza University of Rome
 -- @cite https://doi.org/10.xxxx/yyyyy
 --
 -- @section DEPENDENCIES
 -- - Dependency1: Description or version details.
 -- - Dependency2: Description or version details.
 --
 -- @section LICENSE
 -- This file is part of the Aeneas HyperCompute Platform.
 --
 -- Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 --
 -- @section CHANGELOG
 -- @version 1.0.0-dev - 23th August 2023
 -- - Initial release
 --
 -- @todo
 -- - Complete level vector generator function
 -- - Add training
 --
 -- @see
 -- -
 -- -
 -- -
 --
 --

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity level_vec_gen is
    Port ( level_vec_out : out  STD_LOGIC_VECTOR (63 downto 0);
           frame_index : in  STD_LOGIC_VECTOR (2 downto 0);
           frame_id : in  STD_LOGIC_VECTOR (4 downto 0));
end level_vec_gen;

architecture Behavioral of level_vec_gen is
begin
    process (frame_index, frame_id)
    begin
        -- Update this function to match your requirements
        case frame_index is
            when "000" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0110110011110011111011100000011101101011001100000101111000100011";
                    when "00001" => level_vec_out <= "0111110011110111111011100000011101101011001100000101111000100011";
                    when "00010" => level_vec_out <= "0111110011110111111011100000011101101011001100000101111000100011";
                    when "00011" => level_vec_out <= "0111110011110111111011100000011101101011001100100101111000100011";
                    when "00100" => level_vec_out <= "0111110011110111111011100000011101101011001100100101111000100011";
                    when "00101" => level_vec_out <= "0111110011110111111011100000011101101011001100100101111000100011";
                    when "00110" => level_vec_out <= "0111110011110111111111100000011101101011001100100101111000100011";
                    when "00111" => level_vec_out <= "0111110011110111111111100000011101101011011100100101111000100011";
                    when "01000" => level_vec_out <= "0111110011111111111111100000011101101011011100100101111000100011";
                    when "01001" => level_vec_out <= "0111110011111111111111100000011101101011011100100101111000100011";
                    when "01010" => level_vec_out <= "0111110011111111111111100000011101101011111100100101111001100011";
                    when "01011" => level_vec_out <= "0111111011111111111111100000011101101011111100101101111001100011";
                    when "01100" => level_vec_out <= "0111111011111111111111100000011101101011111100101101111001100011";
                    when "01101" => level_vec_out <= "0111111011111111111111100000011101101011111100101101111001100011";
                    when "01110" => level_vec_out <= "0111111011111111111111100000011101101011111100111101111001100011";
                    when "01111" => level_vec_out <= "0111111011111111111111100000011101101011111100111101111001100011";
                    when "10000" => level_vec_out <= "0111111011111111111111101000011101101011111100111111111001100011";
                    when "10001" => level_vec_out <= "0111111011111111111111101000011111101011111100111111111001100011";
                    when "10010" => level_vec_out <= "0111111011111111111111101000011111101011111100111111111001101011";
                    when "10011" => level_vec_out <= "0111111011111111111111101100011111101011111100111111111011101011";
                    when "10100" => level_vec_out <= "0111111011111111111111101100011111101011111100111111111011111011";
                    when "10101" => level_vec_out <= "0111111011111111111111101100011111101011111100111111111011111011";
                    when "10110" => level_vec_out <= "0111111011111111111111101100011111101011111101111111111011111011";
                    when "10111" => level_vec_out <= "0111111011111111111111101100011111101011111101111111111011111011";
                    when "11000" => level_vec_out <= "0111111011111111111111101100011111111011111101111111111011111011";
                    when "11001" => level_vec_out <= "0111111011111111111111111100011111111011111101111111111111111011";
                    when "11010" => level_vec_out <= "0111111011111111111111111100011111111111111101111111111111111011";
                    when "11011" => level_vec_out <= "1111111011111111111111111110011111111111111101111111111111111011";
                    when "11100" => level_vec_out <= "1111111011111111111111111111011111111111111111111111111111111111";
                    when "11101" => level_vec_out <= "1111111011111111111111111111011111111111111111111111111111111111";
                    when "11110" => level_vec_out <= "1111111011111111111111111111011111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111011111111111111111111111111111111111";
                when others => null;
                end case;
            when "001" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1011001110101111000000000000010001001110000001001011000000101001";
                    when "00001" => level_vec_out <= "1011001110101111000000000000010001001110000001001011100000101001";
                    when "00010" => level_vec_out <= "1011001110101111000000000001010001101110000001001011100000101001";
                    when "00011" => level_vec_out <= "1011001110101111100000000001010001111110000001011011100000101001";
                    when "00100" => level_vec_out <= "1011001110101111100000000001010001111110000001111011100000101001";
                    when "00101" => level_vec_out <= "1011001110101111100100100001010101111110000001111011100000101001";
                    when "00110" => level_vec_out <= "1011001110101111100100100001010101111110000001111011100000101001";
                    when "00111" => level_vec_out <= "1011001110101111100100100001110101111110000101111111100000101001";
                    when "01000" => level_vec_out <= "1011001110101111100100100001110111111110000101111111100000101001";
                    when "01001" => level_vec_out <= "1011001111101111100100100001110111111110001101111111100000101001";
                    when "01010" => level_vec_out <= "1011011111101111100100100001110111111110001101111111100000101001";
                    when "01011" => level_vec_out <= "1011011111101111100100100001110111111110001101111111100000101101";
                    when "01100" => level_vec_out <= "1011011111101111100100100001110111111110001101111111100000101101";
                    when "01101" => level_vec_out <= "1011011111101111100100100001110111111110001101111111101001101101";
                    when "01110" => level_vec_out <= "1011011111101111100100100001110111111110001101111111101001101101";
                    when "01111" => level_vec_out <= "1011011111111111100100100001110111111110001101111111101001101101";
                    when "10000" => level_vec_out <= "1011011111111111100100100011110111111110001101111111101011101101";
                    when "10001" => level_vec_out <= "1011011111111111100100101011110111111110101111111111101011101101";
                    when "10010" => level_vec_out <= "1011011111111111100100101011110111111110111111111111101011101101";
                    when "10011" => level_vec_out <= "1011011111111111110100101011110111111110111111111111101011101101";
                    when "10100" => level_vec_out <= "1011011111111111110100101011110111111110111111111111101111101101";
                    when "10101" => level_vec_out <= "1011111111111111110100111111110111111110111111111111101111101101";
                    when "10110" => level_vec_out <= "1011111111111111110101111111110111111110111111111111101111101111";
                    when "10111" => level_vec_out <= "1111111111111111110101111111110111111110111111111111101111101111";
                    when "11000" => level_vec_out <= "1111111111111111110101111111110111111110111111111111101111101111";
                    when "11001" => level_vec_out <= "1111111111111111110101111111110111111111111111111111101111101111";
                    when "11010" => level_vec_out <= "1111111111111111110101111111110111111111111111111111101111101111";
                    when "11011" => level_vec_out <= "1111111111111111110111111111110111111111111111111111101111101111";
                    when "11100" => level_vec_out <= "1111111111111111110111111111110111111111111111111111101111101111";
                    when "11101" => level_vec_out <= "1111111111111111110111111111110111111111111111111111101111101111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111110111111111111111111111101111101111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111110111111111111111111111111111101111";
                when others => null;
                end case;
            when "010" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1111100000101111101110001110110100110100010110011111101011011010";
                    when "00001" => level_vec_out <= "1111101000101111101110001110110100110100010110011111101011011010";
                    when "00010" => level_vec_out <= "1111101000101111101110001110110100110100010110011111101011011010";
                    when "00011" => level_vec_out <= "1111101000101111101110001110110100110100010110011111101011111010";
                    when "00100" => level_vec_out <= "1111101000101111101110001110110100110100010110011111101011111010";
                    when "00101" => level_vec_out <= "1111101000101111101110001110110110110100010111011111101011111010";
                    when "00110" => level_vec_out <= "1111101001101111101110001110110110110100010111011111101011111110";
                    when "00111" => level_vec_out <= "1111101001101111101110001110110110111100010111011111101011111110";
                    when "01000" => level_vec_out <= "1111101001101111101110011110110110111100010111011111101011111110";
                    when "01001" => level_vec_out <= "1111101001101111101110111110110110111100010111011111101011111110";
                    when "01010" => level_vec_out <= "1111101001111111101111111110110110111100010111011111101011111110";
                    when "01011" => level_vec_out <= "1111101001111111101111111110110110111100010111011111101011111110";
                    when "01100" => level_vec_out <= "1111101101111111101111111110110110111100010111011111101111111110";
                    when "01101" => level_vec_out <= "1111101101111111101111111110110110111100010111011111101111111110";
                    when "01110" => level_vec_out <= "1111101101111111101111111110110110111100010111011111101111111110";
                    when "01111" => level_vec_out <= "1111101101111111101111111110110110111100010111111111101111111110";
                    when "10000" => level_vec_out <= "1111101101111111101111111110110110111100010111111111101111111110";
                    when "10001" => level_vec_out <= "1111101101111111101111111110110110111100010111111111101111111110";
                    when "10010" => level_vec_out <= "1111101101111111101111111110110110111100110111111111101111111110";
                    when "10011" => level_vec_out <= "1111101101111111101111111110110110111100111111111111101111111110";
                    when "10100" => level_vec_out <= "1111101111111111101111111110110110111100111111111111101111111110";
                    when "10101" => level_vec_out <= "1111111111111111101111111110110110111101111111111111101111111110";
                    when "10110" => level_vec_out <= "1111111111111111101111111110110110111111111111111111101111111110";
                    when "10111" => level_vec_out <= "1111111111111111101111111111110110111111111111111111101111111110";
                    when "11000" => level_vec_out <= "1111111111111111101111111111110110111111111111111111101111111110";
                    when "11001" => level_vec_out <= "1111111111111111101111111111110110111111111111111111101111111110";
                    when "11010" => level_vec_out <= "1111111111111111111111111111110111111111111111111111101111111110";
                    when "11011" => level_vec_out <= "1111111111111111111111111111110111111111111111111111101111111110";
                    when "11100" => level_vec_out <= "1111111111111111111111111111110111111111111111111111111111111110";
                    when "11101" => level_vec_out <= "1111111111111111111111111111110111111111111111111111111111111110";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111110";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "011" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1111100100011001001101101111101001101101111000011011110111111001";
                    when "00001" => level_vec_out <= "1111101100011001001101101111101001101101111000011011110111111001";
                    when "00010" => level_vec_out <= "1111101100011001001101101111101001101101111000011011110111111001";
                    when "00011" => level_vec_out <= "1111101100011001001101101111101001101101111000011011110111111001";
                    when "00100" => level_vec_out <= "1111101100011001001101101111101011101101111000011011110111111001";
                    when "00101" => level_vec_out <= "1111101100011001001101101111101011101101111000011011110111111001";
                    when "00110" => level_vec_out <= "1111101100011001001101101111101011101101111000011011110111111001";
                    when "00111" => level_vec_out <= "1111101100011001001101101111101011101101111000011011110111111001";
                    when "01000" => level_vec_out <= "1111101101011001001101101111101011101101111000011011110111111001";
                    when "01001" => level_vec_out <= "1111101101011001001101101111101011101111111000111011111111111001";
                    when "01010" => level_vec_out <= "1111101101011001001101101111101011101111111000111011111111111001";
                    when "01011" => level_vec_out <= "1111101101011001001101101111101011101111111000111011111111111001";
                    when "01100" => level_vec_out <= "1111101101011001001101101111101011101111111000111011111111111001";
                    when "01101" => level_vec_out <= "1111101101011001001101101111101011101111111001111011111111111001";
                    when "01110" => level_vec_out <= "1111101101011001001101101111101011111111111001111011111111111001";
                    when "01111" => level_vec_out <= "1111101101011001001101101111101011111111111001111011111111111001";
                    when "10000" => level_vec_out <= "1111101101011001001101101111101011111111111001111011111111111001";
                    when "10001" => level_vec_out <= "1111101101011001001101101111101111111111111001111011111111111001";
                    when "10010" => level_vec_out <= "1111101101011001001101111111101111111111111001111011111111111001";
                    when "10011" => level_vec_out <= "1111101101011101001101111111101111111111111001111011111111111001";
                    when "10100" => level_vec_out <= "1111101101111101001101111111101111111111111001111011111111111001";
                    when "10101" => level_vec_out <= "1111101101111101001101111111101111111111111001111011111111111001";
                    when "10110" => level_vec_out <= "1111101101111101001101111111101111111111111001111011111111111001";
                    when "10111" => level_vec_out <= "1111101101111101001111111111101111111111111001111011111111111001";
                    when "11000" => level_vec_out <= "1111101101111101001111111111111111111111111001111011111111111101";
                    when "11001" => level_vec_out <= "1111101101111101001111111111111111111111111101111011111111111101";
                    when "11010" => level_vec_out <= "1111101101111101011111111111111111111111111101111011111111111101";
                    when "11011" => level_vec_out <= "1111101101111101011111111111111111111111111101111011111111111101";
                    when "11100" => level_vec_out <= "1111101101111101011111111111111111111111111101111011111111111111";
                    when "11101" => level_vec_out <= "1111111101111101011111111111111111111111111101111111111111111111";
                    when "11110" => level_vec_out <= "1111111111111101011111111111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111101011111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "100" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0111110011111110101011011101010011001001011110110111000001000011";
                    when "00001" => level_vec_out <= "0111110011111110101011011101010011001001011111110111000001000011";
                    when "00010" => level_vec_out <= "0111110011111110101011011101010011001001011111110111000001001011";
                    when "00011" => level_vec_out <= "0111110011111110101011011101010011001001011111110111000001001011";
                    when "00100" => level_vec_out <= "0111110011111110101011011111010011011001011111110111010001001011";
                    when "00101" => level_vec_out <= "0111110011111111101011011111010011011001011111110111010001001011";
                    when "00110" => level_vec_out <= "0111110011111111101011011111010011011001011111110111010001001011";
                    when "00111" => level_vec_out <= "0111110011111111101011011111010011011001011111110111010001001011";
                    when "01000" => level_vec_out <= "0111110011111111101011011111010011011001011111110111010001001011";
                    when "01001" => level_vec_out <= "0111110011111111101011011111010011011001011111110111010001001011";
                    when "01010" => level_vec_out <= "0111110011111111101011011111010011011001011111110111010001001011";
                    when "01011" => level_vec_out <= "0111110011111111111011011111010011011001011111111111010001001011";
                    when "01100" => level_vec_out <= "0111110011111111111011011111010011011001011111111111011001001011";
                    when "01101" => level_vec_out <= "0111110011111111111011011111010011011001011111111111011001001011";
                    when "01110" => level_vec_out <= "0111110011111111111011011111010011011001011111111111011001001011";
                    when "01111" => level_vec_out <= "0111110011111111111011111111010011011001011111111111011001001011";
                    when "10000" => level_vec_out <= "0111110011111111111011111111010011111101011111111111011001001011";
                    when "10001" => level_vec_out <= "0111110111111111111011111111010011111101011111111111011001001011";
                    when "10010" => level_vec_out <= "0111110111111111111011111111010011111101011111111111011001001111";
                    when "10011" => level_vec_out <= "0111110111111111111011111111010011111101011111111111011001001111";
                    when "10100" => level_vec_out <= "0111110111111111111011111111010011111101011111111111011001001111";
                    when "10101" => level_vec_out <= "0111110111111111111011111111011011111111011111111111011001001111";
                    when "10110" => level_vec_out <= "0111110111111111111011111111011011111111011111111111011001001111";
                    when "10111" => level_vec_out <= "0111110111111111111011111111011011111111011111111111011011101111";
                    when "11000" => level_vec_out <= "1111111111111111111011111111111011111111011111111111011011101111";
                    when "11001" => level_vec_out <= "1111111111111111111011111111111011111111011111111111011011101111";
                    when "11010" => level_vec_out <= "1111111111111111111011111111111011111111011111111111011011111111";
                    when "11011" => level_vec_out <= "1111111111111111111011111111111011111111011111111111111111111111";
                    when "11100" => level_vec_out <= "1111111111111111111011111111111011111111011111111111111111111111";
                    when "11101" => level_vec_out <= "1111111111111111111111111111111011111111111111111111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "101" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1001000100000001110110111101010001111000001001100010001000010110";
                    when "00001" => level_vec_out <= "1001000100000001110110111101010001111000001001100010001000010110";
                    when "00010" => level_vec_out <= "1001000100000001110110111101010011111000001001100010001100011110";
                    when "00011" => level_vec_out <= "1001000100000001110110111101010011111000001001100010001100011110";
                    when "00100" => level_vec_out <= "1001000100000001110110111101010011111000001001100010001100011110";
                    when "00101" => level_vec_out <= "1001000100000001110110111101010011111000001001100010001100011111";
                    when "00110" => level_vec_out <= "1001000100000001110110111101010011111000001001101010001100011111";
                    when "00111" => level_vec_out <= "1001000110100001110110111101010011111000001001101010001100011111";
                    when "01000" => level_vec_out <= "1001001110100001110110111101010011111000001001101010001100011111";
                    when "01001" => level_vec_out <= "1001001110100001110110111101010011111000001001101010001100011111";
                    when "01010" => level_vec_out <= "1001001110100001110110111101010011111000001001101010001100011111";
                    when "01011" => level_vec_out <= "1001001110100001110110111111010011111000001001101010001100011111";
                    when "01100" => level_vec_out <= "1101011110100001110110111111010011111000011001111010101100011111";
                    when "01101" => level_vec_out <= "1111011110100001110110111111010111111000011001111010101110011111";
                    when "01110" => level_vec_out <= "1111011110100001110110111111010111111000011001111110101110011111";
                    when "01111" => level_vec_out <= "1111011110100001110111111111010111111000011001111111101110011111";
                    when "10000" => level_vec_out <= "1111011110100001110111111111010111111000011001111111101110011111";
                    when "10001" => level_vec_out <= "1111011110100001110111111111010111111000011001111111101110011111";
                    when "10010" => level_vec_out <= "1111011110100001110111111111010111111000011101111111111110011111";
                    when "10011" => level_vec_out <= "1111011111100101110111111111010111111000011101111111111110011111";
                    when "10100" => level_vec_out <= "1111011111101101110111111111010111111010011101111111111110011111";
                    when "10101" => level_vec_out <= "1111011111101101110111111111011111111010011101111111111110011111";
                    when "10110" => level_vec_out <= "1111011111101101110111111111011111111010011101111111111110011111";
                    when "10111" => level_vec_out <= "1111011111101101110111111111011111111010011101111111111110111111";
                    when "11000" => level_vec_out <= "1111011111101101110111111111011111111010011101111111111110111111";
                    when "11001" => level_vec_out <= "1111011111101111110111111111011111111010011101111111111110111111";
                    when "11010" => level_vec_out <= "1111011111101111110111111111011111111010011101111111111111111111";
                    when "11011" => level_vec_out <= "1111011111101111110111111111011111111010011111111111111111111111";
                    when "11100" => level_vec_out <= "1111111111101111110111111111011111111010011111111111111111111111";
                    when "11101" => level_vec_out <= "1111111111101111110111111111011111111011011111111111111111111111";
                    when "11110" => level_vec_out <= "1111111111101111110111111111011111111011011111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111110111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "110" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0001101000011100100111001010110101101101011110000101010001001000";
                    when "00001" => level_vec_out <= "0001101000011100100111001010110101101101011110000111010001001000";
                    when "00010" => level_vec_out <= "0001101000011100100111001010110101101101011110000111010001001000";
                    when "00011" => level_vec_out <= "0001101000011100110111001011110101101101011110000111010001001000";
                    when "00100" => level_vec_out <= "0001101000011100110111001011110101101101011110000111010001001000";
                    when "00101" => level_vec_out <= "0001101000011100110111001011110101101101011110000111010001001000";
                    when "00110" => level_vec_out <= "0001101001011100110111001011111101111101011110000111010001001000";
                    when "00111" => level_vec_out <= "0001101001011100110111001011111101111101011110100111010001001000";
                    when "01000" => level_vec_out <= "0001101001011100110111001011111111111101011110100111010001001000";
                    when "01001" => level_vec_out <= "0001101001011100110111001011111111111101011110100111010001001000";
                    when "01010" => level_vec_out <= "0001101001011100110111001011111111111101011110100111010001001000";
                    when "01011" => level_vec_out <= "0001101001011100110111001011111111111101011110100111010001001001";
                    when "01100" => level_vec_out <= "0001101001011100110111001011111111111101011110100111010001001001";
                    when "01101" => level_vec_out <= "0001101001011101110111001011111111111101011110100111010001001001";
                    when "01110" => level_vec_out <= "0111101001011101110111001011111111111101011110101111010101001001";
                    when "01111" => level_vec_out <= "0111101001011101110111001011111111111101011110101111010101011001";
                    when "10000" => level_vec_out <= "0111101001011101110111001011111111111101011110111111010101011001";
                    when "10001" => level_vec_out <= "0111101001011101110111011011111111111101011110111111010101011001";
                    when "10010" => level_vec_out <= "0111101001011101110111011011111111111101011110111111010101011001";
                    when "10011" => level_vec_out <= "0111101001011101110111011011111111111101011110111111010101011001";
                    when "10100" => level_vec_out <= "1111101101011101110111011011111111111101011110111111010101011001";
                    when "10101" => level_vec_out <= "1111101101011101110111011011111111111101011110111111010101011001";
                    when "10110" => level_vec_out <= "1111101101011101111111011011111111111101011110111111010111011001";
                    when "10111" => level_vec_out <= "1111111101011101111111011011111111111101011110111111011111011001";
                    when "11000" => level_vec_out <= "1111111101011101111111011011111111111101011110111111011111011001";
                    when "11001" => level_vec_out <= "1111111101011111111111011011111111111101011110111111011111011101";
                    when "11010" => level_vec_out <= "1111111111011111111111011011111111111101011110111111011111011101";
                    when "11011" => level_vec_out <= "1111111111011111111111011111111111111101011110111111011111011101";
                    when "11100" => level_vec_out <= "1111111111011111111111011111111111111101111110111111111111011101";
                    when "11101" => level_vec_out <= "1111111111011111111111011111111111111101111110111111111111111101";
                    when "11110" => level_vec_out <= "1111111111011111111111111111111111111101111110111111111111111111";
                    when "11111" => level_vec_out <= "1111111111011111111111111111111111111111111110111111111111111111";
                when others => null;
                end case;
            when "111" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1100010000101000011100110100100110101100101111101100000100010110";
                    when "00001" => level_vec_out <= "1101010000101000011100110100100110101100101111101100000100010110";
                    when "00010" => level_vec_out <= "1101010000101000011100110100100110101100101111101100100100010111";
                    when "00011" => level_vec_out <= "1101010000101000011100110101100110101100101111101100100100010111";
                    when "00100" => level_vec_out <= "1101011000101000111100110101101110101100101111101100100100010111";
                    when "00101" => level_vec_out <= "1101011000101100111100110101101110101100101111101100100100010111";
                    when "00110" => level_vec_out <= "1101011000101100111100110101101110101100101111101110100100010111";
                    when "00111" => level_vec_out <= "1101011000101100111100110101101110101100101111101110100100010111";
                    when "01000" => level_vec_out <= "1101011000101100111100110101101111101100101111101110101100010111";
                    when "01001" => level_vec_out <= "1101011001101100111100110101101111101100101111111110101100010111";
                    when "01010" => level_vec_out <= "1101011111101100111100110101101111101100101111111111101100010111";
                    when "01011" => level_vec_out <= "1101011111101100111100110101101111101100101111111111101110010111";
                    when "01100" => level_vec_out <= "1101011111101100111100110101101111101100101111111111101110010111";
                    when "01101" => level_vec_out <= "1101011111101101111100110101101111101100101111111111101110010111";
                    when "01110" => level_vec_out <= "1111011111101101111100110101101111101100101111111111101110010111";
                    when "01111" => level_vec_out <= "1111011111101111111100110101101111101100101111111111101110110111";
                    when "10000" => level_vec_out <= "1111011111101111111100110101101111111100101111111111101110110111";
                    when "10001" => level_vec_out <= "1111011111101111111100110101101111111100101111111111101111110111";
                    when "10010" => level_vec_out <= "1111011111101111111100110101101111111100111111111111101111110111";
                    when "10011" => level_vec_out <= "1111011111101111111110110101101111111100111111111111101111110111";
                    when "10100" => level_vec_out <= "1111011111101111111110110101101111111100111111111111101111110111";
                    when "10101" => level_vec_out <= "1111011111101111111110110101101111111100111111111111101111110111";
                    when "10110" => level_vec_out <= "1111111111101111111110110101101111111101111111111111101111110111";
                    when "10111" => level_vec_out <= "1111111111101111111110110101101111111101111111111111101111110111";
                    when "11000" => level_vec_out <= "1111111111101111111110110101111111111101111111111111111111110111";
                    when "11001" => level_vec_out <= "1111111111101111111110110101111111111101111111111111111111111111";
                    when "11010" => level_vec_out <= "1111111111101111111111110101111111111101111111111111111111111111";
                    when "11011" => level_vec_out <= "1111111111111111111111110101111111111101111111111111111111111111";
                    when "11100" => level_vec_out <= "1111111111111111111111110101111111111101111111111111111111111111";
                    when "11101" => level_vec_out <= "1111111111111111111111110111111111111111111111111111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when others => null;
        end case;
    end process;
end Behavioral;