/**
 * @file level_hvec_gen_hdl.hpp
 * @brief This script generates HDL code for generating high-dimensional LEVEL vectors.
 * It is a novel method; for more information, please refer to our paper.
 *
 * @author Saeid Jamili and Marco Angioli
 * @note Author names are listed in alphabetical order.
 * @email <saeid.jamili@uniroma1.it>
 * @email <marco.angioli@uniroma1.it>
 *
 * @contributors
 *
 * @date Created: 24th July 2023
 * @date Last Updated: 23th August 2023
 *
 * @version 1.0.0
 *
 * @institute Sapienza University of Rome
 * @cite https://doi.org/10.xxxx/yyyyy
 *
 * @section DEPENDENCIES
 * - Dependency1: Description or version details.
 * - Dependency2: Description or version details.
 *
 * @section LICENSE
 * This file is part of the Aeneas HyperCompute Platform.
 *
 * Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 *
 * @section CHANGELOG
 * @version 1.0.0-dev - 23th August 2023
 * - Initial release
 *
 * @todo
 * - Complete level vector generator function
 * - Add training
 *
 * @see
 * -
 * -
 * -
 *
 */

module level_hvec_gen #(parameter int DI_PARALLEL_W_BITS = 64) (
  input logic [2:0] frame_index,
  input logic [4:0] frame_id,
  output logic [DI_PARALLEL_W_BITS-1:0] level_vec_out
);
  always_comb begin
    case (frame_index)
      0:
        case (frame_id)
          0:
            level_vec_out = 64'b0110101101101110010010001111000000100111000011010111000001011111;
          1:
            level_vec_out = 64'b0110101101101110010010001111000000100111000011010111001001011111;
          2:
            level_vec_out = 64'b0110101101111110010010011111000010100111000011010111001001011111;
          3:
            level_vec_out = 64'b0110101101111110010010011111000010100111000011010111001001011111;
          4:
            level_vec_out = 64'b0110101101111110010010011111000010100111001011010111001001011111;
          5:
            level_vec_out = 64'b0110101101111110010010011111000010100111101011010111001001011111;
          6:
            level_vec_out = 64'b0110101101111110010010011111000010100111101011010111001001011111;
          7:
            level_vec_out = 64'b0110101101111110010110011111000010100111101011010111101001011111;
          8:
            level_vec_out = 64'b0110101101111110010110011111000010101111101011010111101001011111;
          9:
            level_vec_out = 64'b0110101101111110010110011111000010101111101011010111101001011111;
          10:
            level_vec_out = 64'b0110101101111110010110011111000010101111101011010111101001011111;
          11:
            level_vec_out = 64'b0110101101111110010110011111000010101111101011010111101001111111;
          12:
            level_vec_out = 64'b0110101101111110010110011111000110101111101011010111101001111111;
          13:
            level_vec_out = 64'b0110101101111110010110011111000110101111101011010111101001111111;
          14:
            level_vec_out = 64'b0110101101111110010110011111000110101111101011010111101001111111;
          15:
            level_vec_out = 64'b0110101101111110010110011111010110101111101011010111101001111111;
          16:
            level_vec_out = 64'b0110101101111110110110011111010110101111101111010111101001111111;
          17:
            level_vec_out = 64'b0110101101111110110110011111010110101111101111010111101001111111;
          18:
            level_vec_out = 64'b0110101101111110110110111111010110101111101111010111101001111111;
          19:
            level_vec_out = 64'b0110101101111110110110111111010110101111111111010111101001111111;
          20:
            level_vec_out = 64'b0110101101111110110110111111010110101111111111010111101001111111;
          21:
            level_vec_out = 64'b0111101101111110110110111111010110101111111111010111101001111111;
          22:
            level_vec_out = 64'b0111101111111110110110111111010110101111111111011111101001111111;
          23:
            level_vec_out = 64'b0111101111111110110110111111010110101111111111011111101001111111;
          24:
            level_vec_out = 64'b0111101111111110110110111111011110101111111111111111101001111111;
          25:
            level_vec_out = 64'b0111101111111110111110111111011110101111111111111111101001111111;
          26:
            level_vec_out = 64'b0111101111111110111110111111111110101111111111111111111001111111;
          27:
            level_vec_out = 64'b0111101111111110111110111111111110101111111111111111111101111111;
          28:
            level_vec_out = 64'b1111101111111110111110111111111110101111111111111111111101111111;
          29:
            level_vec_out = 64'b1111111111111110111110111111111111101111111111111111111101111111;
          30:
            level_vec_out = 64'b1111111111111110111110111111111111101111111111111111111101111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111101111111;
        endcase
      1:
        case (frame_id)
          0:
            level_vec_out = 64'b0001110101100101101001011101100100010010001000101000101110010010;
          1:
            level_vec_out = 64'b0001111101100101101001011101100100010110001000101000101110010010;
          2:
            level_vec_out = 64'b0001111101100101101001011101100100010110001000101000101110010010;
          3:
            level_vec_out = 64'b0001111101100101101001011101101100010110001000101000101110010010;
          4:
            level_vec_out = 64'b1001111101100101101001011101101100010110001010101000101110010010;
          5:
            level_vec_out = 64'b1001111101100101101001011101101100010110001010101000101110010010;
          6:
            level_vec_out = 64'b1001111101100101101001011101101100110110001010101100101110010010;
          7:
            level_vec_out = 64'b1001111101100101101001011101101100110110001010101100101110010010;
          8:
            level_vec_out = 64'b1001111101101101101101011101101100110110001010101100111110010010;
          9:
            level_vec_out = 64'b1001111101101101101101011101101101110110101010101100111110010010;
          10:
            level_vec_out = 64'b1001111101101111101101011101101101110111101010101100111110010011;
          11:
            level_vec_out = 64'b1101111101101111101101011101101101110111101010101100111110010011;
          12:
            level_vec_out = 64'b1101111101101111101101011101101101110111111010101100111110010011;
          13:
            level_vec_out = 64'b1101111101101111101101011101101101110111111110101100111110010011;
          14:
            level_vec_out = 64'b1101111111101111101101011101101101110111111110101100111110010011;
          15:
            level_vec_out = 64'b1101111111101111101111011101101101110111111110101100111110010011;
          16:
            level_vec_out = 64'b1101111111101111101111011101101101110111111110101110111110010011;
          17:
            level_vec_out = 64'b1101111111101111101111111111101101110111111110111110111110010011;
          18:
            level_vec_out = 64'b1101111111101111101111111111101111110111111110111110111110010011;
          19:
            level_vec_out = 64'b1101111111101111101111111111101111110111111110111110111110010011;
          20:
            level_vec_out = 64'b1101111111101111101111111111101111110111111110111110111110010011;
          21:
            level_vec_out = 64'b1101111111101111101111111111111111110111111110111110111110010011;
          22:
            level_vec_out = 64'b1101111111101111101111111111111111110111111110111110111110010011;
          23:
            level_vec_out = 64'b1101111111101111101111111111111111110111111110111110111110010011;
          24:
            level_vec_out = 64'b1101111111101111101111111111111111110111111110111110111110110011;
          25:
            level_vec_out = 64'b1101111111101111101111111111111111110111111110111110111110110011;
          26:
            level_vec_out = 64'b1111111111101111101111111111111111110111111110111110111110110011;
          27:
            level_vec_out = 64'b1111111111101111101111111111111111110111111110111110111110110011;
          28:
            level_vec_out = 64'b1111111111101111101111111111111111110111111110111110111110110111;
          29:
            level_vec_out = 64'b1111111111101111101111111111111111110111111110111110111110111111;
          30:
            level_vec_out = 64'b1111111111111111111111111111111111110111111110111111111110111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111110111111111110111111;
        endcase
      2:
        case (frame_id)
          0:
            level_vec_out = 64'b0011011100101000010101110001010001011010100101101001110001110111;
          1:
            level_vec_out = 64'b0011011100101000010101110001010001011010100101101001110001110111;
          2:
            level_vec_out = 64'b0011011100101000010101110001010001011010100101101001110001110111;
          3:
            level_vec_out = 64'b0011011100101000010111110001010001011010100101101001110001110111;
          4:
            level_vec_out = 64'b0011011100101000010111110001010001011010100101101001110001110111;
          5:
            level_vec_out = 64'b0011011100111000010111110001010001011010110101101001110001110111;
          6:
            level_vec_out = 64'b0011011100111000010111110001010001011010110101101001110001110111;
          7:
            level_vec_out = 64'b0011011100111000010111110001010001011010110101101001110001110111;
          8:
            level_vec_out = 64'b0011011100111000010111110001010001011010110101101001110101110111;
          9:
            level_vec_out = 64'b0111011100111000010111110001010001011010110101101001110101110111;
          10:
            level_vec_out = 64'b0111011100111000010111111001010001011010110101101001110101110111;
          11:
            level_vec_out = 64'b0111011100111000010111111001010001011010110101101011110101110111;
          12:
            level_vec_out = 64'b0111011100111000010111111001010001011010110101101011110101110111;
          13:
            level_vec_out = 64'b0111011100111000010111111001010101111010110101101011110101110111;
          14:
            level_vec_out = 64'b0111011100111000010111111001010101111010110111101011110101110111;
          15:
            level_vec_out = 64'b0111011100111000010111111001010101111010110111101011110101110111;
          16:
            level_vec_out = 64'b0111011100111010010111111001010101111010110111101011110101110111;
          17:
            level_vec_out = 64'b0111011110111010010111111001010101111010110111101011110101110111;
          18:
            level_vec_out = 64'b0111011110111010010111111001010101111010110111111011110101110111;
          19:
            level_vec_out = 64'b1111011110111110010111111001110101111010110111111011110101110111;
          20:
            level_vec_out = 64'b1111011110111110011111111001110101111010110111111111111111111111;
          21:
            level_vec_out = 64'b1111011110111110011111111001110101111110110111111111111111111111;
          22:
            level_vec_out = 64'b1111011110111111011111111001110101111110111111111111111111111111;
          23:
            level_vec_out = 64'b1111011110111111011111111001111101111110111111111111111111111111;
          24:
            level_vec_out = 64'b1111111110111111011111111001111101111110111111111111111111111111;
          25:
            level_vec_out = 64'b1111111110111111011111111001111101111110111111111111111111111111;
          26:
            level_vec_out = 64'b1111111110111111011111111001111101111110111111111111111111111111;
          27:
            level_vec_out = 64'b1111111110111111011111111001111101111110111111111111111111111111;
          28:
            level_vec_out = 64'b1111111110111111011111111011111101111110111111111111111111111111;
          29:
            level_vec_out = 64'b1111111110111111011111111011111101111111111111111111111111111111;
          30:
            level_vec_out = 64'b1111111111111111011111111011111111111111111111111111111111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        endcase
      3:
        case (frame_id)
          0:
            level_vec_out = 64'b0101000101100100000100111011101110011011100100101110011010111100;
          1:
            level_vec_out = 64'b0101000101100100000100111011101110011011100100101110011010111100;
          2:
            level_vec_out = 64'b0101000101100100000100111011101110011011101100101110011010111100;
          3:
            level_vec_out = 64'b0101000101100100000100111011101110011011101100101111011010111100;
          4:
            level_vec_out = 64'b0101000101100100010100111011101110011011101100101111011010111100;
          5:
            level_vec_out = 64'b0101001101100100010100111011101110011011101100101111011010111100;
          6:
            level_vec_out = 64'b0111001101100100010100111011101110011011101100101111011010111100;
          7:
            level_vec_out = 64'b0111001101100100010100111011101110011011101100101111011010111100;
          8:
            level_vec_out = 64'b0111001101100100010100111011101110011011101100101111011010111100;
          9:
            level_vec_out = 64'b0111001101100100010100111011101110011011101100101111011010111100;
          10:
            level_vec_out = 64'b0111001101100101010100111011101110011011101100101111011010111100;
          11:
            level_vec_out = 64'b0111001101100101010101111111101110011011101100101111011010111100;
          12:
            level_vec_out = 64'b0111001101100101010101111111111110011011101100101111011010111100;
          13:
            level_vec_out = 64'b0111001101100101010101111111111110011011101100101111011010111100;
          14:
            level_vec_out = 64'b0111001101100101010101111111111110011011101110101111011010111100;
          15:
            level_vec_out = 64'b0111001101100101010101111111111110011011111110101111011010111101;
          16:
            level_vec_out = 64'b0111001101100101010101111111111110011011111110101111011010111101;
          17:
            level_vec_out = 64'b0111001101100101010111111111111110011011111110101111011010111101;
          18:
            level_vec_out = 64'b0111101101100101010111111111111110111011111110101111011010111101;
          19:
            level_vec_out = 64'b0111101101100101010111111111111110111011111110101111011010111111;
          20:
            level_vec_out = 64'b0111101101100101010111111111111110111011111110101111011010111111;
          21:
            level_vec_out = 64'b0111101111100101011111111111111110111011111110101111011010111111;
          22:
            level_vec_out = 64'b0111101111100101011111111111111110111011111110101111011010111111;
          23:
            level_vec_out = 64'b0111101111100101111111111111111110111011111110111111011010111111;
          24:
            level_vec_out = 64'b0111101111101101111111111111111110111011111110111111011010111111;
          25:
            level_vec_out = 64'b0111101111101111111111111111111110111111111110111111011011111111;
          26:
            level_vec_out = 64'b0111101111101111111111111111111110111111111110111111011111111111;
          27:
            level_vec_out = 64'b1111101111101111111111111111111110111111111111111111011111111111;
          28:
            level_vec_out = 64'b1111101111101111111111111111111110111111111111111111011111111111;
          29:
            level_vec_out = 64'b1111101111101111111111111111111110111111111111111111111111111111;
          30:
            level_vec_out = 64'b1111101111101111111111111111111110111111111111111111111111111111;
          31:
            level_vec_out = 64'b1111101111101111111111111111111110111111111111111111111111111111;
        endcase
      4:
        case (frame_id)
          0:
            level_vec_out = 64'b0111000010101010011111110011010001110100110000100111101011100010;
          1:
            level_vec_out = 64'b1111001010101010011111110011010001110100110000100111101011100010;
          2:
            level_vec_out = 64'b1111001010101010011111110011010001110100110010100111101011100010;
          3:
            level_vec_out = 64'b1111001010111010011111110011010001110100110010100111111011100010;
          4:
            level_vec_out = 64'b1111001010111011011111110011010001110100110010101111111011100010;
          5:
            level_vec_out = 64'b1111001010111011011111110011010001110100110010101111111011100010;
          6:
            level_vec_out = 64'b1111001010111011011111110011010001110100111011101111111011100010;
          7:
            level_vec_out = 64'b1111001010111011011111110111010001110100111011101111111011101010;
          8:
            level_vec_out = 64'b1111001010111011011111110111010001110100111011101111111011101010;
          9:
            level_vec_out = 64'b1111001010111011011111110111010001110101111011101111111011101010;
          10:
            level_vec_out = 64'b1111101010111011011111110111010001110101111011101111111011101010;
          11:
            level_vec_out = 64'b1111101010111011011111110111010001110101111011101111111011101010;
          12:
            level_vec_out = 64'b1111101010111011011111110111010101110101111111101111111011101010;
          13:
            level_vec_out = 64'b1111101010111011011111110111010101110101111111101111111011101010;
          14:
            level_vec_out = 64'b1111101010111011011111110111110101110101111111101111111011101010;
          15:
            level_vec_out = 64'b1111101010111011011111110111111101110101111111101111111011101010;
          16:
            level_vec_out = 64'b1111101010111011011111110111111101110101111111101111111011101010;
          17:
            level_vec_out = 64'b1111101010111011011111110111111101110101111111101111111011101010;
          18:
            level_vec_out = 64'b1111101010111011011111110111111101110101111111101111111011101010;
          19:
            level_vec_out = 64'b1111101010111011011111110111111101110101111111101111111011101010;
          20:
            level_vec_out = 64'b1111101010111111011111110111111101110101111111101111111011101010;
          21:
            level_vec_out = 64'b1111101010111111011111110111111101110101111111101111111011101010;
          22:
            level_vec_out = 64'b1111101010111111011111111111111101111101111111101111111011101010;
          23:
            level_vec_out = 64'b1111101010111111011111111111111101111101111111101111111111101010;
          24:
            level_vec_out = 64'b1111101011111111011111111111111101111111111111101111111111101010;
          25:
            level_vec_out = 64'b1111101011111111011111111111111101111111111111101111111111101011;
          26:
            level_vec_out = 64'b1111111011111111111111111111111101111111111111101111111111101011;
          27:
            level_vec_out = 64'b1111111011111111111111111111111101111111111111101111111111101011;
          28:
            level_vec_out = 64'b1111111111111111111111111111111101111111111111101111111111101111;
          29:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111101111111111101111;
          30:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111101111111111101111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        endcase
      5:
        case (frame_id)
          0:
            level_vec_out = 64'b0010101110000101000110110100010001010101000011001001100011010101;
          1:
            level_vec_out = 64'b0010101110000101000110110100010001011101000011001001100011010101;
          2:
            level_vec_out = 64'b0010101110000101000110110100010001011101000011001011100011010101;
          3:
            level_vec_out = 64'b0010101110100101000110110100010001011101000011001011100011010101;
          4:
            level_vec_out = 64'b0010101110100101000110110100010001011101000011001011100011010101;
          5:
            level_vec_out = 64'b0010101110100101000110110100010001011101000011001011100011010101;
          6:
            level_vec_out = 64'b1010101110100101000110110110010001011101000011001011100011010101;
          7:
            level_vec_out = 64'b1010101110100101000110110110010001011101000011001011100011010101;
          8:
            level_vec_out = 64'b1010101110110101000110110110010001011101000011001011100011010101;
          9:
            level_vec_out = 64'b1010101110110101000110110110010001011101000011001111100011110101;
          10:
            level_vec_out = 64'b1010101110110101000110110110111001011101000011001111100011110101;
          11:
            level_vec_out = 64'b1010101110110101000110110110111001111101000011001111100011110101;
          12:
            level_vec_out = 64'b1010101110110101000110111110111001111101000011001111100011110101;
          13:
            level_vec_out = 64'b1010101110110101000110111110111101111101001011001111100011110101;
          14:
            level_vec_out = 64'b1010101110110101000110111110111101111101001011001111100011110101;
          15:
            level_vec_out = 64'b1010101110110101000110111110111101111101001011101111100011110101;
          16:
            level_vec_out = 64'b1010101110110101000110111110111101111111001011101111100111110101;
          17:
            level_vec_out = 64'b1010101110110101000110111110111101111111011011101111100111110101;
          18:
            level_vec_out = 64'b1010101110110101001110111110111101111111011011101111110111110101;
          19:
            level_vec_out = 64'b1010101110110101001111111111111101111111011011101111110111110101;
          20:
            level_vec_out = 64'b1010101110110101001111111111111101111111011011101111110111110101;
          21:
            level_vec_out = 64'b1010101110110101001111111111111101111111011011101111110111111101;
          22:
            level_vec_out = 64'b1010101110110101001111111111111101111111011011101111110111111101;
          23:
            level_vec_out = 64'b1011111110110101001111111111111101111111011011101111110111111101;
          24:
            level_vec_out = 64'b1011111110110101001111111111111101111111011011101111110111111101;
          25:
            level_vec_out = 64'b1011111111110101001111111111111101111111011011101111110111111101;
          26:
            level_vec_out = 64'b1011111111110101001111111111111111111111011011101111110111111101;
          27:
            level_vec_out = 64'b1011111111110101001111111111111111111111011111101111111111111111;
          28:
            level_vec_out = 64'b1011111111111101001111111111111111111111111111101111111111111111;
          29:
            level_vec_out = 64'b1111111111111101001111111111111111111111111111101111111111111111;
          30:
            level_vec_out = 64'b1111111111111101011111111111111111111111111111111111111111111111;
          31:
            level_vec_out = 64'b1111111111111101011111111111111111111111111111111111111111111111;
        endcase
      6:
        case (frame_id)
          0:
            level_vec_out = 64'b1001001011101000010111101100100110110100011100000001101001001010;
          1:
            level_vec_out = 64'b1001001011101000010111111100100110110101011100000001101001001010;
          2:
            level_vec_out = 64'b1001001011101000010111111100110110110101011100000001101001001010;
          3:
            level_vec_out = 64'b1001001011101000010111111100110110110101011100000001101001001010;
          4:
            level_vec_out = 64'b1001001011111000010111111100110110110101011100000001101001001010;
          5:
            level_vec_out = 64'b1001101011111000010111111111110110110101011100000001101001001010;
          6:
            level_vec_out = 64'b1001101011111000010111111111110110110111011100000001101001001010;
          7:
            level_vec_out = 64'b1001101111111000010111111111110110110111111100000001101001001010;
          8:
            level_vec_out = 64'b1001101111111000011111111111110110110111111101000001101001001010;
          9:
            level_vec_out = 64'b1001101111111000011111111111110110110111111101000001101001001010;
          10:
            level_vec_out = 64'b1001101111111000011111111111110110110111111101000001101001001010;
          11:
            level_vec_out = 64'b1001101111111010011111111111110110110111111101000101101001001010;
          12:
            level_vec_out = 64'b1001101111111010011111111111110110110111111101000101101001101010;
          13:
            level_vec_out = 64'b1011101111111110011111111111110110110111111101010101101001101010;
          14:
            level_vec_out = 64'b1011101111111110111111111111110110110111111101010101101001101010;
          15:
            level_vec_out = 64'b1011111111111110111111111111110110110111111101010101101001111010;
          16:
            level_vec_out = 64'b1011111111111111111111111111110110110111111101010101101001111010;
          17:
            level_vec_out = 64'b1011111111111111111111111111110110110111111101110101101001111010;
          18:
            level_vec_out = 64'b1011111111111111111111111111110110110111111101110101101001111010;
          19:
            level_vec_out = 64'b1011111111111111111111111111110110110111111101110101101101111010;
          20:
            level_vec_out = 64'b1111111111111111111111111111110110110111111101110101101111111010;
          21:
            level_vec_out = 64'b1111111111111111111111111111110110110111111101110101111111111010;
          22:
            level_vec_out = 64'b1111111111111111111111111111110110110111111101110111111111111110;
          23:
            level_vec_out = 64'b1111111111111111111111111111110110111111111111110111111111111110;
          24:
            level_vec_out = 64'b1111111111111111111111111111110110111111111111110111111111111110;
          25:
            level_vec_out = 64'b1111111111111111111111111111110110111111111111110111111111111110;
          26:
            level_vec_out = 64'b1111111111111111111111111111110110111111111111110111111111111110;
          27:
            level_vec_out = 64'b1111111111111111111111111111110110111111111111110111111111111111;
          28:
            level_vec_out = 64'b1111111111111111111111111111111110111111111111110111111111111111;
          29:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111110111111111111111;
          30:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        endcase
      7:
        case (frame_id)
          0:
            level_vec_out = 64'b1111100110110111011110001010101110111101101011011010110110001111;
          1:
            level_vec_out = 64'b1111100110110111011110001010101110111101101011011010110110001111;
          2:
            level_vec_out = 64'b1111100110110111011110001010101110111101101011011110110110001111;
          3:
            level_vec_out = 64'b1111101110110111011111001010101110111101101011011110110110001111;
          4:
            level_vec_out = 64'b1111101110110111011111001010101110111101101011011111110110001111;
          5:
            level_vec_out = 64'b1111101110110111011111001010101111111101101011011111110110001111;
          6:
            level_vec_out = 64'b1111101110110111011111001010101111111101101011011111110110001111;
          7:
            level_vec_out = 64'b1111101110110111011111001010101111111101101111111111110110001111;
          8:
            level_vec_out = 64'b1111101110110111011111001010101111111101101111111111110110001111;
          9:
            level_vec_out = 64'b1111111110110111111111001010101111111101101111111111110110001111;
          10:
            level_vec_out = 64'b1111111110110111111111001010101111111101101111111111110110001111;
          11:
            level_vec_out = 64'b1111111110110111111111001010101111111101101111111111110110001111;
          12:
            level_vec_out = 64'b1111111110110111111111001011101111111101101111111111110110001111;
          13:
            level_vec_out = 64'b1111111110110111111111001011101111111101101111111111110110001111;
          14:
            level_vec_out = 64'b1111111110110111111111001011101111111111101111111111110111011111;
          15:
            level_vec_out = 64'b1111111110110111111111001011101111111111101111111111110111011111;
          16:
            level_vec_out = 64'b1111111110110111111111101011101111111111101111111111110111011111;
          17:
            level_vec_out = 64'b1111111110110111111111111011101111111111101111111111110111011111;
          18:
            level_vec_out = 64'b1111111110110111111111111011101111111111101111111111111111011111;
          19:
            level_vec_out = 64'b1111111110110111111111111011101111111111101111111111111111011111;
          20:
            level_vec_out = 64'b1111111110110111111111111011101111111111101111111111111111011111;
          21:
            level_vec_out = 64'b1111111110110111111111111011101111111111101111111111111111111111;
          22:
            level_vec_out = 64'b1111111110110111111111111011101111111111101111111111111111111111;
          23:
            level_vec_out = 64'b1111111110110111111111111011101111111111101111111111111111111111;
          24:
            level_vec_out = 64'b1111111110110111111111111111101111111111101111111111111111111111;
          25:
            level_vec_out = 64'b1111111111111111111111111111101111111111101111111111111111111111;
          26:
            level_vec_out = 64'b1111111111111111111111111111101111111111111111111111111111111111;
          27:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
          28:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
          29:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
          30:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        endcase
    endcase
  end
endmodule