----
 -- @file level_hvec_gen_hdl.hpp
 -- @brief This script generates HDL code for generating high-dimensional LEVEL vectors.
 -- It is a novel method; for more information, please refer to our paper.
 --
 -- @author Saeid Jamili and Marco Angioli
 -- @note Author names are listed in alphabetical order.
 -- @email <saeid.jamili@uniroma1.it>
 -- @email <marco.angioli@uniroma1.it>
 --
 -- @contributors
 --
 -- @date Created: 24th July 2023
 -- @date Last Updated: 23th August 2023
 --
 -- @version 1.0.0
 --
 -- @institute Sapienza University of Rome
 -- @cite https://doi.org/10.xxxx/yyyyy
 --
 -- @section DEPENDENCIES
 -- - Dependency1: Description or version details.
 -- - Dependency2: Description or version details.
 --
 -- @section LICENSE
 -- This file is part of the Aeneas HyperCompute Platform.
 --
 -- Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 --
 -- @section CHANGELOG
 -- @version 1.0.0-dev - 23th August 2023
 -- - Initial release
 --
 -- @todo
 -- - Complete level vector generator function
 -- - Add training
 --
 -- @see
 -- -
 -- -
 -- -
 --
 --

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity level_vec_gen is
    Port ( level_vec_out : out  STD_LOGIC_VECTOR (63 downto 0);
           frame_index : in  STD_LOGIC_VECTOR (2 downto 0);
           frame_id : in  STD_LOGIC_VECTOR (4 downto 0));
end level_vec_gen;

architecture Behavioral of level_vec_gen is
begin
    process (frame_index, frame_id)
    begin
        -- Update this function to match your requirements
        case frame_index is
            when "000" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1110010100010001000010111001100101010000011000000101100100101110";
                    when "00001" => level_vec_out <= "1110010110010001000010111001100101011000011000000101100100101110";
                    when "00010" => level_vec_out <= "1110010111010011000010111001100101011000011000000101100100101110";
                    when "00011" => level_vec_out <= "1110010111010011000010111001100101011000011000000101100100101110";
                    when "00100" => level_vec_out <= "1110010111010011000010111001100101011000011000100101100100101110";
                    when "00101" => level_vec_out <= "1110010111010011000010111001100101011000011000100101100100101110";
                    when "00110" => level_vec_out <= "1110010111010011000010111001101101011000011000100101100100111110";
                    when "00111" => level_vec_out <= "1110010111011011000010111001101111011000011000100101100100111110";
                    when "01000" => level_vec_out <= "1110010111011011000010111001101111011000011000100101100100111110";
                    when "01001" => level_vec_out <= "1110010111011011000010111001111111011000011000100101100100111110";
                    when "01010" => level_vec_out <= "1110010111011011000010111001111111011000011000100101100100111110";
                    when "01011" => level_vec_out <= "1110010111011011000010111001111111011000011000100101100100111110";
                    when "01100" => level_vec_out <= "1110010111011011100010111001111111011001011010100101100100111110";
                    when "01101" => level_vec_out <= "1110011111011011100010111011111111011001011010100101100100111110";
                    when "01110" => level_vec_out <= "1111011111011011100010111011111111011001111111100111100100111110";
                    when "01111" => level_vec_out <= "1111011111011011101010111011111111111001111111100111100100111110";
                    when "10000" => level_vec_out <= "1111011111011011101010111011111111111001111111100111100100111110";
                    when "10001" => level_vec_out <= "1111011111011011111010111011111111111001111111100111100101111110";
                    when "10010" => level_vec_out <= "1111011111011111111010111011111111111001111111101111100111111110";
                    when "10011" => level_vec_out <= "1111011111011111111110111011111111111001111111101111100111111110";
                    when "10100" => level_vec_out <= "1111011111011111111110111111111111111011111111101111110111111110";
                    when "10101" => level_vec_out <= "1111011111011111111111111111111111111011111111101111110111111110";
                    when "10110" => level_vec_out <= "1111011111011111111111111111111111111011111111101111110111111110";
                    when "10111" => level_vec_out <= "1111011111011111111111111111111111111011111111101111110111111110";
                    when "11000" => level_vec_out <= "1111011111011111111111111111111111111011111111101111110111111110";
                    when "11001" => level_vec_out <= "1111011111011111111111111111111111111011111111101111110111111110";
                    when "11010" => level_vec_out <= "1111011111011111111111111111111111111011111111101111110111111110";
                    when "11011" => level_vec_out <= "1111011111011111111111111111111111111011111111101111110111111110";
                    when "11100" => level_vec_out <= "1111011111011111111111111111111111111011111111101111110111111111";
                    when "11101" => level_vec_out <= "1111011111011111111111111111111111111111111111101111110111111111";
                    when "11110" => level_vec_out <= "1111111111011111111111111111111111111111111111101111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111101111111111111111";
                when others => null;
                end case;
            when "001" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0010110111110111011111001100111101111010110011101101000110000100";
                    when "00001" => level_vec_out <= "1010110111110111011111001100111101111010110011101101000110000100";
                    when "00010" => level_vec_out <= "1010110111110111011111001100111101111010110011101101000110000100";
                    when "00011" => level_vec_out <= "1010110111110111011111001100111101111010110011101101000110000100";
                    when "00100" => level_vec_out <= "1010110111110111011111001100111101111010110011101101000110000100";
                    when "00101" => level_vec_out <= "1010110111110111011111001100111101111010110011111101000110000100";
                    when "00110" => level_vec_out <= "1010110111110111011111001100111111111010110011111101000110000100";
                    when "00111" => level_vec_out <= "1010110111110111011111001100111111111010110011111101000110000100";
                    when "01000" => level_vec_out <= "1010110111110111011111001100111111111010110111111101100110001100";
                    when "01001" => level_vec_out <= "1010110111110111011111001100111111111010110111111101100110001100";
                    when "01010" => level_vec_out <= "1010110111110111011111001110111111111010110111111101100110001100";
                    when "01011" => level_vec_out <= "1010110111110111011111001110111111111110110111111101100110001100";
                    when "01100" => level_vec_out <= "1010110111110111011111001110111111111110110111111101100110001100";
                    when "01101" => level_vec_out <= "1010110111110111011111001110111111111110110111111101100110001100";
                    when "01110" => level_vec_out <= "1010110111110111011111001110111111111110110111111101100110001100";
                    when "01111" => level_vec_out <= "1010110111110111011111011110111111111110110111111101100110001100";
                    when "10000" => level_vec_out <= "1010110111110111011111011110111111111110110111111101100110001100";
                    when "10001" => level_vec_out <= "1110110111110111011111111110111111111110110111111101100110001110";
                    when "10010" => level_vec_out <= "1110110111110111011111111110111111111110110111111101100110001110";
                    when "10011" => level_vec_out <= "1110110111110111011111111110111111111110110111111101100110011110";
                    when "10100" => level_vec_out <= "1110110111110111011111111110111111111110110111111101100110011110";
                    when "10101" => level_vec_out <= "1110110111110111011111111110111111111111110111111101100110011110";
                    when "10110" => level_vec_out <= "1110110111110111011111111110111111111111110111111101100110011111";
                    when "10111" => level_vec_out <= "1110110111111111011111111110111111111111110111111101100110011111";
                    when "11000" => level_vec_out <= "1110110111111111111111111110111111111111111111111101100110011111";
                    when "11001" => level_vec_out <= "1111110111111111111111111110111111111111111111111101110110011111";
                    when "11010" => level_vec_out <= "1111110111111111111111111110111111111111111111111101110110111111";
                    when "11011" => level_vec_out <= "1111110111111111111111111110111111111111111111111101110111111111";
                    when "11100" => level_vec_out <= "1111110111111111111111111110111111111111111111111101110111111111";
                    when "11101" => level_vec_out <= "1111110111111111111111111110111111111111111111111101110111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111110111111111111111111111101110111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111101110111111111";
                when others => null;
                end case;
            when "010" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1000111101110111010000010011000001010110110000101101000001100010";
                    when "00001" => level_vec_out <= "1000111101110111010000010011000001010110110000101101001001100010";
                    when "00010" => level_vec_out <= "1000111101110111010000010011100001010110110000101101001001100010";
                    when "00011" => level_vec_out <= "1000111101110111010000010011100001110110110000101101101001100010";
                    when "00100" => level_vec_out <= "1000111101110111010000010011100001110110110000101101101001100010";
                    when "00101" => level_vec_out <= "1000111101110111010000010011100001110110110001101101101001100010";
                    when "00110" => level_vec_out <= "1000111101110111110010010011100011110110110001101101101001100010";
                    when "00111" => level_vec_out <= "1000111101110111110010010011100011110110110001101101101001100010";
                    when "01000" => level_vec_out <= "1000111101110111110010010011101011110110110011101101101001100010";
                    when "01001" => level_vec_out <= "1000111101110111110010010011101011110110110011101101101001100010";
                    when "01010" => level_vec_out <= "1000111101110111110010010011101011110110110011101101101001100010";
                    when "01011" => level_vec_out <= "1000111101110111110010010011101011110110110011101101101001100010";
                    when "01100" => level_vec_out <= "1000111101110111110010010111101011111110110011101101101001100010";
                    when "01101" => level_vec_out <= "1000111101110111111010010111101011111110110011101101101001100010";
                    when "01110" => level_vec_out <= "1000111101110111111010010111101011111110110111101101101001100010";
                    when "01111" => level_vec_out <= "1000111101110111111010010111101011111110110111101101101011100010";
                    when "10000" => level_vec_out <= "1000111101110111111010010111101011111110110111101101101011100010";
                    when "10001" => level_vec_out <= "1000111101110111111010010111101011111110110111101101101011100010";
                    when "10010" => level_vec_out <= "1000111111110111111010010111101011111110110111101101101011100010";
                    when "10011" => level_vec_out <= "1000111111110111111010010111101111111110110111101101101111100010";
                    when "10100" => level_vec_out <= "1001111111110111111110110111101111111110110111101101101111100010";
                    when "10101" => level_vec_out <= "1001111111110111111110111111101111111110110111101101101111100011";
                    when "10110" => level_vec_out <= "1001111111111111111110111111101111111110110111111101101111100011";
                    when "10111" => level_vec_out <= "1001111111111111111110111111101111111110110111111101101111100011";
                    when "11000" => level_vec_out <= "1001111111111111111110111111101111111110110111111101101111100011";
                    when "11001" => level_vec_out <= "1001111111111111111110111111101111111110110111111101101111101111";
                    when "11010" => level_vec_out <= "1101111111111111111111111111101111111110110111111101101111101111";
                    when "11011" => level_vec_out <= "1101111111111111111111111111101111111111110111111101101111101111";
                    when "11100" => level_vec_out <= "1101111111111111111111111111101111111111111111111101111111111111";
                    when "11101" => level_vec_out <= "1111111111111111111111111111111111111111111111111101111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "011" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1101000111010111010100100011110011010010001001100001000111111110";
                    when "00001" => level_vec_out <= "1101000111010111010100110011110011010010001001100001000111111110";
                    when "00010" => level_vec_out <= "1101000111010111010100110011110011010010001001100001000111111110";
                    when "00011" => level_vec_out <= "1101000111010111010100110011110011010010001001100011000111111110";
                    when "00100" => level_vec_out <= "1101000111010111010100110011110011010010001001100011000111111110";
                    when "00101" => level_vec_out <= "1101101111010111010110110011110011010010001011100011000111111110";
                    when "00110" => level_vec_out <= "1101101111010111010110110011110011010010001011100011000111111110";
                    when "00111" => level_vec_out <= "1101101111010111010110110111110011010010001011100011000111111110";
                    when "01000" => level_vec_out <= "1101101111010111010110110111110011010010001011100011000111111110";
                    when "01001" => level_vec_out <= "1101101111010111010110111111110011010010001011100011000111111111";
                    when "01010" => level_vec_out <= "1101111111010111010110111111110011010010001011100011000111111111";
                    when "01011" => level_vec_out <= "1101111111010111010110111111110011010010001011100011000111111111";
                    when "01100" => level_vec_out <= "1101111111010111010110111111110011010010001011100011000111111111";
                    when "01101" => level_vec_out <= "1101111111010111010110111111110011010010011011100011100111111111";
                    when "01110" => level_vec_out <= "1101111111010111010110111111110011010010011011100011100111111111";
                    when "01111" => level_vec_out <= "1101111111010111010110111111110011010010111011100111100111111111";
                    when "10000" => level_vec_out <= "1101111111010111010110111111110011010011111011100111101111111111";
                    when "10001" => level_vec_out <= "1101111111010111010111111111110011010011111011100111101111111111";
                    when "10010" => level_vec_out <= "1101111111010111010111111111110011011011111011100111101111111111";
                    when "10011" => level_vec_out <= "1101111111010111010111111111110011011011111111100111101111111111";
                    when "10100" => level_vec_out <= "1101111111010111010111111111110011011011111111100111101111111111";
                    when "10101" => level_vec_out <= "1101111111010111010111111111110011011011111111100111101111111111";
                    when "10110" => level_vec_out <= "1101111111111111110111111111110011011011111111100111101111111111";
                    when "10111" => level_vec_out <= "1101111111111111110111111111110011011011111111100111101111111111";
                    when "11000" => level_vec_out <= "1101111111111111110111111111110011011011111111100111101111111111";
                    when "11001" => level_vec_out <= "1101111111111111110111111111110011011011111111100111101111111111";
                    when "11010" => level_vec_out <= "1101111111111111110111111111110011011111111111100111101111111111";
                    when "11011" => level_vec_out <= "1101111111111111110111111111110011011111111111110111101111111111";
                    when "11100" => level_vec_out <= "1101111111111111110111111111110011111111111111110111101111111111";
                    when "11101" => level_vec_out <= "1111111111111111111111111111110011111111111111110111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111110111111111111111110111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111110111111111111111111111111111111111";
                when others => null;
                end case;
            when "100" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1001010010101000101101001011011101110001111111100011000001001111";
                    when "00001" => level_vec_out <= "1001010010101000101101001011011101110001111111100011000001001111";
                    when "00010" => level_vec_out <= "1001010110101000101101001011011101110001111111100011000001001111";
                    when "00011" => level_vec_out <= "1001010110101000101101001011011101110001111111100011000001001111";
                    when "00100" => level_vec_out <= "1001010110101000101101001011011101110001111111100011000001001111";
                    when "00101" => level_vec_out <= "1001010110101000101101001011011101110001111111100011000001011111";
                    when "00110" => level_vec_out <= "1001010110101000101111001011011101110001111111100011000001011111";
                    when "00111" => level_vec_out <= "1001010110101000101111001011011101111001111111100011000001011111";
                    when "01000" => level_vec_out <= "1001010110101000101111001011011101111001111111100011000001111111";
                    when "01001" => level_vec_out <= "1001010110101000101111001011011101111001111111101011000001111111";
                    when "01010" => level_vec_out <= "1001011110101001101111001011011101111001111111101011000001111111";
                    when "01011" => level_vec_out <= "1001011110101001101111001011011101111001111111101011000001111111";
                    when "01100" => level_vec_out <= "1001011110101001101111001011011101111001111111101011000001111111";
                    when "01101" => level_vec_out <= "1001011110101001101111001011011101111001111111101111000001111111";
                    when "01110" => level_vec_out <= "1101011110101001101111001111011101111001111111101111000001111111";
                    when "01111" => level_vec_out <= "1111011110101001111111001111011101111001111111101111000001111111";
                    when "10000" => level_vec_out <= "1111011110101111111111001111011101111001111111101111000001111111";
                    when "10001" => level_vec_out <= "1111011110101111111111001111011101111001111111101111000001111111";
                    when "10010" => level_vec_out <= "1111011110101111111111001111011101111001111111101111000001111111";
                    when "10011" => level_vec_out <= "1111111110101111111111001111011101111011111111101111000011111111";
                    when "10100" => level_vec_out <= "1111111110101111111111001111011101111011111111101111000011111111";
                    when "10101" => level_vec_out <= "1111111110101111111111101111011101111011111111101111000011111111";
                    when "10110" => level_vec_out <= "1111111110101111111111101111011101111011111111101111000011111111";
                    when "10111" => level_vec_out <= "1111111110101111111111101111011101111011111111111111000011111111";
                    when "11000" => level_vec_out <= "1111111110101111111111101111011101111111111111111111000111111111";
                    when "11001" => level_vec_out <= "1111111110101111111111101111011101111111111111111111000111111111";
                    when "11010" => level_vec_out <= "1111111110101111111111101111111101111111111111111111100111111111";
                    when "11011" => level_vec_out <= "1111111110101111111111101111111101111111111111111111101111111111";
                    when "11100" => level_vec_out <= "1111111110101111111111101111111101111111111111111111101111111111";
                    when "11101" => level_vec_out <= "1111111110101111111111101111111101111111111111111111101111111111";
                    when "11110" => level_vec_out <= "1111111111101111111111101111111101111111111111111111101111111111";
                    when "11111" => level_vec_out <= "1111111111101111111111101111111101111111111111111111111111111111";
                when others => null;
                end case;
            when "101" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0011011101011000000001110100100101111110111011110101001100101011";
                    when "00001" => level_vec_out <= "0011011101011000000001110100100101111110111011110101001110101011";
                    when "00010" => level_vec_out <= "0011011101011001000001110101100101111110111011110101001110101011";
                    when "00011" => level_vec_out <= "0111011101011101000001110111100101111110111011110101001110101011";
                    when "00100" => level_vec_out <= "0111011101011101000001110111100101111110111011110101001110101011";
                    when "00101" => level_vec_out <= "0111011101011111000001110111100101111110111011110101001110101011";
                    when "00110" => level_vec_out <= "0111011101011111000001110111100101111110111011110101001110101011";
                    when "00111" => level_vec_out <= "0111011101011111000001110111101101111110111011110101001110101011";
                    when "01000" => level_vec_out <= "0111011111011111000001110111101101111110111011110101001110101011";
                    when "01001" => level_vec_out <= "0111011111011111000001110111101101111110111011110101001110101011";
                    when "01010" => level_vec_out <= "0111011111011111000001110111101101111110111011110101001110111011";
                    when "01011" => level_vec_out <= "0111011111011111000001110111101101111110111011110101011110111011";
                    when "01100" => level_vec_out <= "0111011111011111010001110111101101111110111011110101011110111011";
                    when "01101" => level_vec_out <= "0111011111011111010001110111101101111110111011110101011111111011";
                    when "01110" => level_vec_out <= "0111011111011111010001110111101101111110111011110101011111111011";
                    when "01111" => level_vec_out <= "0111011111011111010001110111101101111110111011110101011111111011";
                    when "10000" => level_vec_out <= "1111011111011111010001110111101101111110111011110101011111111011";
                    when "10001" => level_vec_out <= "1111011111011111010001110111101101111110111011110101111111111011";
                    when "10010" => level_vec_out <= "1111011111011111010001110111101101111110111011110101111111111011";
                    when "10011" => level_vec_out <= "1111011111011111010001110111101101111110111011110101111111111011";
                    when "10100" => level_vec_out <= "1111011111011111011001110111101101111110111011110101111111111011";
                    when "10101" => level_vec_out <= "1111011111111111011001110111101101111110111011110101111111111011";
                    when "10110" => level_vec_out <= "1111011111111111011101110111101101111110111011110101111111111011";
                    when "10111" => level_vec_out <= "1111111111111111011101111111101101111110111011110101111111111111";
                    when "11000" => level_vec_out <= "1111111111111111011101111111101111111110111011111101111111111111";
                    when "11001" => level_vec_out <= "1111111111111111011101111111111111111111111111111101111111111111";
                    when "11010" => level_vec_out <= "1111111111111111011101111111111111111111111111111101111111111111";
                    when "11011" => level_vec_out <= "1111111111111111011101111111111111111111111111111101111111111111";
                    when "11100" => level_vec_out <= "1111111111111111011101111111111111111111111111111101111111111111";
                    when "11101" => level_vec_out <= "1111111111111111111111111111111111111111111111111101111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111111111111101111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111101111111111111";
                when others => null;
                end case;
            when "110" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1111011001001111011100001111010001011101011111000100110010010110";
                    when "00001" => level_vec_out <= "1111011001001111011100001111010001011101011111000100110010010110";
                    when "00010" => level_vec_out <= "1111011001001111011101001111010001011101011111000100110010110110";
                    when "00011" => level_vec_out <= "1111011001001111011101001111010001011101011111000100110010110110";
                    when "00100" => level_vec_out <= "1111011011001111011101001111010011011101011111010100111010110110";
                    when "00101" => level_vec_out <= "1111011011001111011101001111010011011101011111010100111010110110";
                    when "00110" => level_vec_out <= "1111011011001111011111001111010011011101011111010100111010110110";
                    when "00111" => level_vec_out <= "1111011011001111011111001111010011111101011111010100111010110110";
                    when "01000" => level_vec_out <= "1111011011001111011111001111010011111101011111010101111010110110";
                    when "01001" => level_vec_out <= "1111011011101111011111001111110011111101011111010101111010110110";
                    when "01010" => level_vec_out <= "1111011011101111011111001111110011111101011111010111111010110110";
                    when "01011" => level_vec_out <= "1111011011101111111111011111111111111101011111010111111010110110";
                    when "01100" => level_vec_out <= "1111011011101111111111011111111111111101011111010111111010110110";
                    when "01101" => level_vec_out <= "1111011011111111111111011111111111111101011111010111111010110110";
                    when "01110" => level_vec_out <= "1111011011111111111111011111111111111101011111010111111010110110";
                    when "01111" => level_vec_out <= "1111011011111111111111011111111111111101011111010111111010110110";
                    when "10000" => level_vec_out <= "1111011011111111111111011111111111111101011111010111111010111110";
                    when "10001" => level_vec_out <= "1111011011111111111111011111111111111101111111010111111010111110";
                    when "10010" => level_vec_out <= "1111111011111111111111011111111111111101111111010111111010111110";
                    when "10011" => level_vec_out <= "1111111011111111111111011111111111111101111111010111111010111110";
                    when "10100" => level_vec_out <= "1111111011111111111111011111111111111101111111010111111010111110";
                    when "10101" => level_vec_out <= "1111111011111111111111111111111111111101111111010111111010111110";
                    when "10110" => level_vec_out <= "1111111011111111111111111111111111111111111111010111111010111110";
                    when "10111" => level_vec_out <= "1111111011111111111111111111111111111111111111010111111011111110";
                    when "11000" => level_vec_out <= "1111111011111111111111111111111111111111111111010111111011111110";
                    when "11001" => level_vec_out <= "1111111011111111111111111111111111111111111111010111111111111110";
                    when "11010" => level_vec_out <= "1111111011111111111111111111111111111111111111010111111111111110";
                    when "11011" => level_vec_out <= "1111111011111111111111111111111111111111111111010111111111111111";
                    when "11100" => level_vec_out <= "1111111011111111111111111111111111111111111111010111111111111111";
                    when "11101" => level_vec_out <= "1111111011111111111111111111111111111111111111010111111111111111";
                    when "11110" => level_vec_out <= "1111111011111111111111111111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "111" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0011110001010011100011001100100001000111000110000001000000101111";
                    when "00001" => level_vec_out <= "0011110001011011100011001100100001100111000110000001000000101111";
                    when "00010" => level_vec_out <= "0011110001011011100011001100100001100111000110000001000000101111";
                    when "00011" => level_vec_out <= "0011110001011011100011001110100001101111000110000001000000101111";
                    when "00100" => level_vec_out <= "0011110001111011110011001110100001101111000110000101000000101111";
                    when "00101" => level_vec_out <= "0011110001111011110011001110100001101111000110000101000000101111";
                    when "00110" => level_vec_out <= "0011110001111011110011001110100001101111000110000101000000101111";
                    when "00111" => level_vec_out <= "0011110001111011110011001110100001101111000111010101000000101111";
                    when "01000" => level_vec_out <= "0011110001111011110011001110100001101111000111010101000000101111";
                    when "01001" => level_vec_out <= "0111110101111011110011001110100001101111000111010101000000101111";
                    when "01010" => level_vec_out <= "0111110101111011110011001110100011101111000111010101000100101111";
                    when "01011" => level_vec_out <= "0111110101111011110011101110100011101111000111010101000110101111";
                    when "01100" => level_vec_out <= "0111110101111011111011111110100011101111000111010101000110101111";
                    when "01101" => level_vec_out <= "0111110101111011111011111110100011101111000111010101000110101111";
                    when "01110" => level_vec_out <= "0111110101111011111011111110100011101111000111010101000110101111";
                    when "01111" => level_vec_out <= "0111110101111011111011111110100011101111000111010101000110101111";
                    when "10000" => level_vec_out <= "0111110101111011111011111110101011101111100111010101000110101111";
                    when "10001" => level_vec_out <= "0111110101111011111011111110101011101111100111010101000110101111";
                    when "10010" => level_vec_out <= "0111111101111011111011111110101011101111100111110101000110101111";
                    when "10011" => level_vec_out <= "0111111101111011111011111110101011101111100111110101000110101111";
                    when "10100" => level_vec_out <= "0111111101111111111011111110101011101111100111110101000110101111";
                    when "10101" => level_vec_out <= "0111111101111111111011111110101011101111100111110101000110111111";
                    when "10110" => level_vec_out <= "0111111101111111111011111110101011101111100111110101000110111111";
                    when "10111" => level_vec_out <= "1111111101111111111011111110101011101111100111110101010110111111";
                    when "11000" => level_vec_out <= "1111111111111111111011111110111011101111100111110101010110111111";
                    when "11001" => level_vec_out <= "1111111111111111111011111110111011101111100111110101010110111111";
                    when "11010" => level_vec_out <= "1111111111111111111011111110111011101111101111110101011110111111";
                    when "11011" => level_vec_out <= "1111111111111111111011111111111011111111101111111101011110111111";
                    when "11100" => level_vec_out <= "1111111111111111111011111111111111111111101111111111111110111111";
                    when "11101" => level_vec_out <= "1111111111111111111011111111111111111111101111111111111110111111";
                    when "11110" => level_vec_out <= "1111111111111111111011111111111111111111101111111111111110111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when others => null;
        end case;
    end process;
end Behavioral;