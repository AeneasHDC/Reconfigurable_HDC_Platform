/**
 * @file level_hvec_gen_hdl.hpp
 * @brief This script generates HDL code for generating high-dimensional LEVEL vectors.
 * It is a novel method; for more information, please refer to our paper.
 *
 * @author Saeid Jamili and Marco Angioli
 * @note Author names are listed in alphabetical order.
 * @email <saeid.jamili@uniroma1.it>
 * @email <marco.angioli@uniroma1.it>
 *
 * @contributors
 *
 * @date Created: 24th July 2023
 * @date Last Updated: 23th August 2023
 *
 * @version 1.0.0
 *
 * @institute Sapienza University of Rome
 * @cite https://doi.org/10.xxxx/yyyyy
 *
 * @section DEPENDENCIES
 * - Dependency1: Description or version details.
 * - Dependency2: Description or version details.
 *
 * @section LICENSE
 * This file is part of the Aeneas HyperCompute Platform.
 *
 * Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 *
 * @section CHANGELOG
 * @version 1.0.0-dev - 23th August 2023
 * - Initial release
 *
 * @todo
 * - Complete level vector generator function
 * - Add training
 *
 * @see
 * -
 * -
 * -
 *
 */

module level_hvec_gen #(parameter int DI_PARALLEL_W_BITS = 64) (
  input logic [2:0] frame_index,
  input logic [4:0] frame_id,
  output logic [DI_PARALLEL_W_BITS-1:0] level_vec_out
);
  always_comb begin
    case (frame_index)
      0:
        case (frame_id)
          0:
            level_vec_out = 64'b0010000110011001001100000000111011001110110010001010010100100010;
          1:
            level_vec_out = 64'b0010000110011001001100000000111011001110110010001010010100100010;
          2:
            level_vec_out = 64'b0010000110011001001100010000111011001110110010001010010100100010;
          3:
            level_vec_out = 64'b0010000110011001001100010000111011001110110010001010010100100010;
          4:
            level_vec_out = 64'b0010001110011001001100010000111011001110110010001010010100100110;
          5:
            level_vec_out = 64'b0010001110011001001100010000111011001110110010001011010100100110;
          6:
            level_vec_out = 64'b1010001110011001001110010000111011001110110010001011010100100110;
          7:
            level_vec_out = 64'b1010001110011001001110010000111011001110111010001011010100100110;
          8:
            level_vec_out = 64'b1010001110011001001110010000111011001110111010011011010100100110;
          9:
            level_vec_out = 64'b1010001110011001011110010000111011001110111010011011010100100110;
          10:
            level_vec_out = 64'b1010001110011001111111010000111011001110111010011011010100100110;
          11:
            level_vec_out = 64'b1010001110011001111111010000111011001110111010011011010100100110;
          12:
            level_vec_out = 64'b1011001110011001111111011000111011001110111010011011010100100110;
          13:
            level_vec_out = 64'b1011001110011001111111011000111011001110111010011011010100100110;
          14:
            level_vec_out = 64'b1011001110011001111111011000111011001110111010011011010100100110;
          15:
            level_vec_out = 64'b1011001110011001111111011000111011001110111010011011010100100110;
          16:
            level_vec_out = 64'b1011101110011001111111011000111011001110111010011011010100100110;
          17:
            level_vec_out = 64'b1011101110111001111111011000111011101110111010011011010100100110;
          18:
            level_vec_out = 64'b1111101110111001111111011000111011101110111010011011010110100110;
          19:
            level_vec_out = 64'b1111101110111001111111111000111011101110111010011011010110100110;
          20:
            level_vec_out = 64'b1111111110111001111111111000111011101111111010011011010110100110;
          21:
            level_vec_out = 64'b1111111111111001111111111000111011111111111010011011010110100111;
          22:
            level_vec_out = 64'b1111111111111001111111111000111011111111111010011011010110100111;
          23:
            level_vec_out = 64'b1111111111111001111111111000111011111111111010011011010110101111;
          24:
            level_vec_out = 64'b1111111111111001111111111010111111111111111010011011010110101111;
          25:
            level_vec_out = 64'b1111111111111101111111111010111111111111111010011011110110101111;
          26:
            level_vec_out = 64'b1111111111111101111111111010111111111111111010011011110110101111;
          27:
            level_vec_out = 64'b1111111111111101111111111010111111111111111111011011110110101111;
          28:
            level_vec_out = 64'b1111111111111101111111111011111111111111111111011011110110101111;
          29:
            level_vec_out = 64'b1111111111111101111111111111111111111111111111111011110110101111;
          30:
            level_vec_out = 64'b1111111111111101111111111111111111111111111111111111110110101111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111110101111;
        endcase
      1:
        case (frame_id)
          0:
            level_vec_out = 64'b0111111111110110011111010010111110101111101110010010000110011011;
          1:
            level_vec_out = 64'b1111111111110110011111010010111110101111101110010010000110011011;
          2:
            level_vec_out = 64'b1111111111110110111111010010111110101111101110011010100110011011;
          3:
            level_vec_out = 64'b1111111111110110111111010010111110101111101110011010100110011011;
          4:
            level_vec_out = 64'b1111111111110110111111010010111110101111101110011010100110011011;
          5:
            level_vec_out = 64'b1111111111110110111111010010111110101111101110011011100110011111;
          6:
            level_vec_out = 64'b1111111111110110111111010010111110101111101111011011110110011111;
          7:
            level_vec_out = 64'b1111111111110110111111010010111110101111101111011011110110011111;
          8:
            level_vec_out = 64'b1111111111110110111111010010111110101111101111011011110110011111;
          9:
            level_vec_out = 64'b1111111111110110111111010010111110101111101111011011110110011111;
          10:
            level_vec_out = 64'b1111111111110110111111010010111110101111101111011011110110011111;
          11:
            level_vec_out = 64'b1111111111110110111111010010111110101111101111011011110110011111;
          12:
            level_vec_out = 64'b1111111111110110111111010010111110101111101111011011110110011111;
          13:
            level_vec_out = 64'b1111111111110110111111010010111110101111101111011011110110011111;
          14:
            level_vec_out = 64'b1111111111110110111111010010111110101111101111011011111110011111;
          15:
            level_vec_out = 64'b1111111111110110111111010011111111101111101111011011111110011111;
          16:
            level_vec_out = 64'b1111111111110110111111010011111111101111101111011011111110011111;
          17:
            level_vec_out = 64'b1111111111110110111111010011111111111111101111011011111110111111;
          18:
            level_vec_out = 64'b1111111111110110111111010011111111111111101111011111111110111111;
          19:
            level_vec_out = 64'b1111111111110110111111110011111111111111101111011111111110111111;
          20:
            level_vec_out = 64'b1111111111110110111111110011111111111111101111011111111110111111;
          21:
            level_vec_out = 64'b1111111111110110111111110011111111111111101111011111111110111111;
          22:
            level_vec_out = 64'b1111111111110110111111110011111111111111101111011111111110111111;
          23:
            level_vec_out = 64'b1111111111110110111111110011111111111111101111011111111110111111;
          24:
            level_vec_out = 64'b1111111111110110111111111011111111111111101111011111111110111111;
          25:
            level_vec_out = 64'b1111111111110111111111111011111111111111101111011111111111111111;
          26:
            level_vec_out = 64'b1111111111110111111111111011111111111111101111011111111111111111;
          27:
            level_vec_out = 64'b1111111111110111111111111111111111111111111111011111111111111111;
          28:
            level_vec_out = 64'b1111111111110111111111111111111111111111111111011111111111111111;
          29:
            level_vec_out = 64'b1111111111110111111111111111111111111111111111011111111111111111;
          30:
            level_vec_out = 64'b1111111111110111111111111111111111111111111111111111111111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        endcase
      2:
        case (frame_id)
          0:
            level_vec_out = 64'b0011101111100110100010011110100101010101110010100111100001110010;
          1:
            level_vec_out = 64'b0011101111100110100011011111100111010101110010100111100001110010;
          2:
            level_vec_out = 64'b0011101111100110100011011111100111010101110010100111100001110010;
          3:
            level_vec_out = 64'b0011101111101110100011011111100111011101110010100111100001110010;
          4:
            level_vec_out = 64'b0011101111101110100011011111100111011101110010100111100001110010;
          5:
            level_vec_out = 64'b0011101111101110100011011111100111011101110010100111100001110010;
          6:
            level_vec_out = 64'b0011101111101110110011011111100111011101110010100111100001110010;
          7:
            level_vec_out = 64'b0011101111101110110011011111100111011101110010100111100101110011;
          8:
            level_vec_out = 64'b0011101111101110110011011111101111011101110010100111110101110011;
          9:
            level_vec_out = 64'b0011101111101110110011011111101111011101111010100111110101110011;
          10:
            level_vec_out = 64'b0011101111101110110011111111101111011101111010100111110101110011;
          11:
            level_vec_out = 64'b0011101111101110110011111111101111011101111011100111110101110011;
          12:
            level_vec_out = 64'b0011101111101110110011111111111111011101111011100111110101110011;
          13:
            level_vec_out = 64'b0111101111101110111011111111111111011101111011100111110101110011;
          14:
            level_vec_out = 64'b0111101111101110111011111111111111011101111011100111110101110011;
          15:
            level_vec_out = 64'b0111101111101110111011111111111111011101111011100111110101110011;
          16:
            level_vec_out = 64'b0111101111101111111011111111111111011101111011110111110101110011;
          17:
            level_vec_out = 64'b0111101111101111111011111111111111011101111011110111110101110011;
          18:
            level_vec_out = 64'b0111111111101111111011111111111111011101111011110111110101110011;
          19:
            level_vec_out = 64'b0111111111101111111011111111111111011101111011110111110101110011;
          20:
            level_vec_out = 64'b0111111111101111111011111111111111011101111011110111110101110011;
          21:
            level_vec_out = 64'b0111111111101111111011111111111111011101111011110111110101110111;
          22:
            level_vec_out = 64'b0111111111101111111111111111111111011101111011110111110111110111;
          23:
            level_vec_out = 64'b1111111111101111111111111111111111011101111111110111110111111111;
          24:
            level_vec_out = 64'b1111111111101111111111111111111111011101111111110111110111111111;
          25:
            level_vec_out = 64'b1111111111101111111111111111111111011101111111110111110111111111;
          26:
            level_vec_out = 64'b1111111111101111111111111111111111011101111111110111110111111111;
          27:
            level_vec_out = 64'b1111111111101111111111111111111111011101111111110111110111111111;
          28:
            level_vec_out = 64'b1111111111111111111111111111111111011101111111110111110111111111;
          29:
            level_vec_out = 64'b1111111111111111111111111111111111011101111111111111111111111111;
          30:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        endcase
      3:
        case (frame_id)
          0:
            level_vec_out = 64'b0001100101101100000010111000011111001000011011110011100100000100;
          1:
            level_vec_out = 64'b0001100101101100000010111000011111001000011011110011100100000100;
          2:
            level_vec_out = 64'b0001100101101100000010111000011111001000011011110011100100000100;
          3:
            level_vec_out = 64'b0001100101101100000010111010011111001000011011110011100100000100;
          4:
            level_vec_out = 64'b0001100101101100000110111010011111001010011011110011100100000100;
          5:
            level_vec_out = 64'b0001100101111100000110111010011111101010011011110011100100000100;
          6:
            level_vec_out = 64'b0001100101111100000110111010011111101010011011110011100100000100;
          7:
            level_vec_out = 64'b0001100101111110000110111010011111101110111011110011100100000100;
          8:
            level_vec_out = 64'b0001101101111110000110111010011111111110111011110011100100000100;
          9:
            level_vec_out = 64'b0011101101111110000110111010011111111110111011110011100100000100;
          10:
            level_vec_out = 64'b0011101101111110000110111010011111111111111011110011100101000100;
          11:
            level_vec_out = 64'b0011101101111110000110111010011111111111111011110011100101000100;
          12:
            level_vec_out = 64'b0011101101111110000110111010011111111111111011110011110101000100;
          13:
            level_vec_out = 64'b0011101101111110000110111010011111111111111011110011110101000100;
          14:
            level_vec_out = 64'b0011101101111110000110111110011111111111111011110011110101010100;
          15:
            level_vec_out = 64'b1011101101111110000110111110111111111111111011110011110101010100;
          16:
            level_vec_out = 64'b1011101101111110000110111110111111111111111011110011110101010100;
          17:
            level_vec_out = 64'b1011101101111110000110111110111111111111111011111011110101010101;
          18:
            level_vec_out = 64'b1011101111111110000110111110111111111111111011111011110101010101;
          19:
            level_vec_out = 64'b1011101111111110100110111110111111111111111011111111110101010111;
          20:
            level_vec_out = 64'b1011101111111110100110111110111111111111111011111111111101010111;
          21:
            level_vec_out = 64'b1011101111111110100110111110111111111111111011111111111101010111;
          22:
            level_vec_out = 64'b1011101111111110100110111110111111111111111011111111111101010111;
          23:
            level_vec_out = 64'b1011101111111110101110111110111111111111111011111111111101010111;
          24:
            level_vec_out = 64'b1011101111111110101110111110111111111111111011111111111101010111;
          25:
            level_vec_out = 64'b1011101111111110101110111110111111111111111011111111111101010111;
          26:
            level_vec_out = 64'b1011111111111110101111111110111111111111111011111111111101010111;
          27:
            level_vec_out = 64'b1011111111111110111111111110111111111111111011111111111101010111;
          28:
            level_vec_out = 64'b1011111111111110111111111110111111111111111011111111111111010111;
          29:
            level_vec_out = 64'b1011111111111110111111111110111111111111111011111111111111110111;
          30:
            level_vec_out = 64'b1011111111111110111111111111111111111111111011111111111111110111;
          31:
            level_vec_out = 64'b1011111111111110111111111111111111111111111011111111111111111111;
        endcase
      4:
        case (frame_id)
          0:
            level_vec_out = 64'b0110010100011010000100010001110011011010101110110011110100001001;
          1:
            level_vec_out = 64'b0110010100011010000100010001110011011010101110110011110100001001;
          2:
            level_vec_out = 64'b0110010100011010000100010001110011011010101110110011110100001001;
          3:
            level_vec_out = 64'b0110010100011010000100010001110011011010101110110011110100001001;
          4:
            level_vec_out = 64'b0110010110011110000100010001111011011010101110110011110100001001;
          5:
            level_vec_out = 64'b0110010110011110000100010001111111011010101110110011110100001001;
          6:
            level_vec_out = 64'b0110010110011110000100010001111111011010101110110011110100001001;
          7:
            level_vec_out = 64'b0111010110011110000100010001111111011010101110110011110100001001;
          8:
            level_vec_out = 64'b0111010110011110000100010001111111011110101110110011110100001001;
          9:
            level_vec_out = 64'b0111010110011110000100010001111111011110111110110011110100001001;
          10:
            level_vec_out = 64'b0111010110011110000100010001111111011110111110110011110100001001;
          11:
            level_vec_out = 64'b0111010110011110000100010001111111011110111110110011110100001001;
          12:
            level_vec_out = 64'b0111010110011110000101010001111111011110111110110011110100001001;
          13:
            level_vec_out = 64'b0111010110011110000111110001111111011110111110110011110100001001;
          14:
            level_vec_out = 64'b0111010110011110000111110001111111011110111110110011110110001001;
          15:
            level_vec_out = 64'b0111010110111110000111110001111111011110111110110011110110001011;
          16:
            level_vec_out = 64'b0111010110111110010111110011111111011110111111110011110110001011;
          17:
            level_vec_out = 64'b0111010110111110010111110011111111011110111111110011110110001011;
          18:
            level_vec_out = 64'b0111010110111110010111110011111111011110111111110011110110001011;
          19:
            level_vec_out = 64'b0111010110111110010111110011111111011110111111111011110110001011;
          20:
            level_vec_out = 64'b0111011110111110010111110011111111011110111111111011111110001011;
          21:
            level_vec_out = 64'b0111111110111110010111110011111111011110111111111011111110001011;
          22:
            level_vec_out = 64'b0111111111111110110111110111111111011110111111111111111110001111;
          23:
            level_vec_out = 64'b0111111111111110110111110111111111011110111111111111111110001111;
          24:
            level_vec_out = 64'b0111111111111110110111110111111111011110111111111111111110001111;
          25:
            level_vec_out = 64'b0111111111111110111111110111111111011110111111111111111110001111;
          26:
            level_vec_out = 64'b0111111111111110111111110111111111011110111111111111111110111111;
          27:
            level_vec_out = 64'b1111111111111110111111110111111111011110111111111111111110111111;
          28:
            level_vec_out = 64'b1111111111111110111111110111111111011111111111111111111110111111;
          29:
            level_vec_out = 64'b1111111111111110111111111111111111011111111111111111111110111111;
          30:
            level_vec_out = 64'b1111111111111110111111111111111111011111111111111111111111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111011111111111111111111111111111;
        endcase
      5:
        case (frame_id)
          0:
            level_vec_out = 64'b1101000010011100101101110101110000100010010001101000110011101011;
          1:
            level_vec_out = 64'b1101000010011100111101110101110000100110010001101000110011101011;
          2:
            level_vec_out = 64'b1101000011011100111101110101110001110110010001101000110011101011;
          3:
            level_vec_out = 64'b1101000011011101111101110101110001110110110001101000110011101011;
          4:
            level_vec_out = 64'b1101000011011101111101110101110001110110110101101000110011101011;
          5:
            level_vec_out = 64'b1101000011011101111101111101110001110110110101101000110011101011;
          6:
            level_vec_out = 64'b1101000011011101111101111101110001110110110101101000110011101011;
          7:
            level_vec_out = 64'b1101000011011101111101111101110001110110110101101000110011101011;
          8:
            level_vec_out = 64'b1101000011011101111101111101110001110110110101101000110011111011;
          9:
            level_vec_out = 64'b1101100011011101111101111101110001110110110101101000110011111011;
          10:
            level_vec_out = 64'b1101100011011101111101111101110001111110110101101000110011111011;
          11:
            level_vec_out = 64'b1101100011011101111111111101110001111110110101101000110011111011;
          12:
            level_vec_out = 64'b1101100011011101111111111111110001111110110101101010110011111011;
          13:
            level_vec_out = 64'b1101100011011101111111111111110001111110110101101010110011111111;
          14:
            level_vec_out = 64'b1101100011011101111111111111110011111110110101101010110011111111;
          15:
            level_vec_out = 64'b1101100011011111111111111111110011111110110101101010110011111111;
          16:
            level_vec_out = 64'b1101100011011111111111111111110011111110110101101010110011111111;
          17:
            level_vec_out = 64'b1101100011011111111111111111110011111110110101101010110011111111;
          18:
            level_vec_out = 64'b1101110011011111111111111111110011111110110111101010110011111111;
          19:
            level_vec_out = 64'b1101110011111111111111111111110011111110110111101010110011111111;
          20:
            level_vec_out = 64'b1101110011111111111111111111110011111110110111101010110011111111;
          21:
            level_vec_out = 64'b1101110011111111111111111111110011111110110111101110110011111111;
          22:
            level_vec_out = 64'b1101110011111111111111111111110011111110110111101110110011111111;
          23:
            level_vec_out = 64'b1101110011111111111111111111110011111110111111101110110011111111;
          24:
            level_vec_out = 64'b1101110011111111111111111111110111111111111111101111110011111111;
          25:
            level_vec_out = 64'b1101110011111111111111111111110111111111111111101111110111111111;
          26:
            level_vec_out = 64'b1101110011111111111111111111111111111111111111101111110111111111;
          27:
            level_vec_out = 64'b1101110011111111111111111111111111111111111111101111110111111111;
          28:
            level_vec_out = 64'b1111110011111111111111111111111111111111111111101111110111111111;
          29:
            level_vec_out = 64'b1111110011111111111111111111111111111111111111111111110111111111;
          30:
            level_vec_out = 64'b1111111011111111111111111111111111111111111111111111110111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111110111111111;
        endcase
      6:
        case (frame_id)
          0:
            level_vec_out = 64'b0110101001111100110011101011100111001010011001011100001001010000;
          1:
            level_vec_out = 64'b0110101001111100110011101011100111011010011001011100001001010000;
          2:
            level_vec_out = 64'b0110101011111100110011101011100111011010011001011100001001010000;
          3:
            level_vec_out = 64'b0110101011111110110011101011100111011010011001011100001001010000;
          4:
            level_vec_out = 64'b0110101011111110110011101011100111011010011001011100001001010000;
          5:
            level_vec_out = 64'b0110101011111110110011101011100111011010011001011100001001010000;
          6:
            level_vec_out = 64'b0110101011111110110011101011100111011010011001111100001001010100;
          7:
            level_vec_out = 64'b0110101011111110110011101011100111011010011001111100001001010100;
          8:
            level_vec_out = 64'b0110101011111110110011101011100111011010011001111100001001010100;
          9:
            level_vec_out = 64'b0110101011111110110011101011101111011110011001111100001001010100;
          10:
            level_vec_out = 64'b0110101011111110110011101011101111011110011001111100001001010100;
          11:
            level_vec_out = 64'b0110111011111110110011101011101111011110011001111100101011010100;
          12:
            level_vec_out = 64'b0110111011111110110011101011101111011110011001111100101011010100;
          13:
            level_vec_out = 64'b0110111011111110110011111011101111111110011001111100101011010100;
          14:
            level_vec_out = 64'b0110111011111110110011111011101111111110011001111100101111010100;
          15:
            level_vec_out = 64'b0110111011111110110011111011101111111110011001111100101111010101;
          16:
            level_vec_out = 64'b0110111011111110111011111011101111111110011001111100101111010101;
          17:
            level_vec_out = 64'b0110111011111110111011111011101111111110111001111101101111010101;
          18:
            level_vec_out = 64'b0110111011111110111011111011101111111110111001111101101111010101;
          19:
            level_vec_out = 64'b0110111011111110111011111011101111111110111001111101101111010101;
          20:
            level_vec_out = 64'b0110111011111110111011111011101111111110111001111101101111010101;
          21:
            level_vec_out = 64'b0110111011111110111111111011101111111110111001111101101111010101;
          22:
            level_vec_out = 64'b0110111011111110111111111011111111111110111001111101101111010101;
          23:
            level_vec_out = 64'b0110111011111110111111111011111111111110111001111101101111010111;
          24:
            level_vec_out = 64'b0110111011111110111111111011111111111110111101111101101111010111;
          25:
            level_vec_out = 64'b0110111011111110111111111011111111111110111101111111101111010111;
          26:
            level_vec_out = 64'b0110111111111110111111111011111111111110111111111111101111010111;
          27:
            level_vec_out = 64'b0110111111111110111111111011111111111110111111111111101111110111;
          28:
            level_vec_out = 64'b1110111111111110111111111111111111111110111111111111111111110111;
          29:
            level_vec_out = 64'b1110111111111110111111111111111111111110111111111111111111111111;
          30:
            level_vec_out = 64'b1110111111111111111111111111111111111110111111111111111111111111;
          31:
            level_vec_out = 64'b1110111111111111111111111111111111111111111111111111111111111111;
        endcase
      7:
        case (frame_id)
          0:
            level_vec_out = 64'b0011100110010111000111100100010100011101010100111001011110110101;
          1:
            level_vec_out = 64'b0011100110010111000111100100010100011101010100111001011110111101;
          2:
            level_vec_out = 64'b0011100110010111000111100100010100011101010100111001011110111101;
          3:
            level_vec_out = 64'b0011100110010111000111100100010100011101010100111011011111111101;
          4:
            level_vec_out = 64'b0011100110010111000111100100010100011101010100111011011111111101;
          5:
            level_vec_out = 64'b1011100110010111000111100100010100011101010100111011011111111101;
          6:
            level_vec_out = 64'b1011100110010111000111100100010110011101010100111011011111111101;
          7:
            level_vec_out = 64'b1011100110010111000111100100010110011101010110111011011111111101;
          8:
            level_vec_out = 64'b1011100110010111000111100100010110011101010110111111011111111101;
          9:
            level_vec_out = 64'b1011100110010111000111100100010110011101010111111111011111111101;
          10:
            level_vec_out = 64'b1011100110010111100111100100010110011101010111111111011111111111;
          11:
            level_vec_out = 64'b1011111110010111100111101100010110011101010111111111011111111111;
          12:
            level_vec_out = 64'b1011111110010111100111101100110110011101010111111111011111111111;
          13:
            level_vec_out = 64'b1011111110010111100111101101110110011101010111111111011111111111;
          14:
            level_vec_out = 64'b1011111110010111100111101101111110011101011111111111011111111111;
          15:
            level_vec_out = 64'b1011111110010111100111101101111110011101011111111111011111111111;
          16:
            level_vec_out = 64'b1011111110011111100111101101111110011101011111111111011111111111;
          17:
            level_vec_out = 64'b1011111110011111100111101101111110011101011111111111011111111111;
          18:
            level_vec_out = 64'b1011111111011111100111101101111110011101011111111111011111111111;
          19:
            level_vec_out = 64'b1011111111011111101111101101111110011101011111111111011111111111;
          20:
            level_vec_out = 64'b1011111111011111111111101111111110011111011111111111011111111111;
          21:
            level_vec_out = 64'b1011111111011111111111101111111110011111011111111111111111111111;
          22:
            level_vec_out = 64'b1011111111011111111111101111111110011111011111111111111111111111;
          23:
            level_vec_out = 64'b1011111111011111111111101111111110111111011111111111111111111111;
          24:
            level_vec_out = 64'b1111111111011111111111101111111110111111011111111111111111111111;
          25:
            level_vec_out = 64'b1111111111011111111111101111111111111111011111111111111111111111;
          26:
            level_vec_out = 64'b1111111111011111111111101111111111111111111111111111111111111111;
          27:
            level_vec_out = 64'b1111111111111111111111101111111111111111111111111111111111111111;
          28:
            level_vec_out = 64'b1111111111111111111111101111111111111111111111111111111111111111;
          29:
            level_vec_out = 64'b1111111111111111111111101111111111111111111111111111111111111111;
          30:
            level_vec_out = 64'b1111111111111111111111101111111111111111111111111111111111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        endcase
    endcase
  end
endmodule