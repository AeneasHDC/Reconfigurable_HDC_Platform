-- Configuration file for VHDL
constant VERBOS_DISABLE : string := 0;
constant VERBOS_L1 : string := 1;
constant VERBOS_L2 : string := 2;
constant VERBOS : string := VERBOS_L1;
constant WINDOWS : string := 0;
constant LINUX : string := 1;
constant MAC : string := 2;
constant OS : string := WINDOWS;
constant FPGA : string := 0;
constant MICROCONTROLER : string := 1;
constant SOFT_PROCESSOR : string := 2;
constant DEVICE_TYPE : string := FPGA;
constant description : string := "Conversion Modes and Configurations";
constant TARGET_DEVICE : string := "xczu9eg-ffvb1156-2-e";
constant AMD_ZYBO : string := 0;
constant AMD_ZEDBOARD : string := 1;
constant AMD_ZCU106 : string := 2;
constant AMD_ZCU102 : string := 3;
constant AMD_VCU108 : string := 4;
constant TARGET_BOARD : string := AMD_ZCU102;
constant OP_FREQ : string := 20;
constant USE_VIV_EN : string := 1;
constant VIV_OPT_DEFAULT : string := 0;
constant VIV_OPT_RESOURCE : string := 1;
constant VIV_OPT_SPEED : string := 2;
constant VIV_OPT_PERFORMANCE : string := 3;
constant VIV_OPT_METHOD : string := VIV_OPT_DEFAULT;
constant HLS : string := 0;
constant SYSTEM_VERILOG : string := 1;
constant VHDL : string := 2;
constant VERILOG : string := 3;
constant HDL_LANG : string := HLS;
constant PYTHON : string := 4;
constant MATLAB : string := 5;
constant CPP : string := 6;
constant C : string := 7;
constant RUST : string := 8;
constant MODEL_LANG : string := PYTHON;
constant DS_NAME : string := "EMG";
constant DS_SIZE : string := 186036;
constant DS_TRAIN_SIZE : string := 372106;
constant DS_TEST_SIZE : string := 148830;
constant DS_VALIDATION_SIZE : string := 372106;
constant DS_FEATURE_SIZE : string := 4;
constant DS_DATA_TYPE : string := "FP";
constant DS_DATA_RANGE_MIN : string := 0;
constant DS_DATA_RANGE_MAX : string := 21;
constant DS_CLASSES_SIZE : string := 5;
constant TRAIN_ON_HW : string := 0;
constant RETRAIN_ON_HW : string := 0;
constant EPOCH : string := 10;
constant HD_DIM : string := 256;
constant BINARY : string := 0;
constant BIPOLAR : string := 1;
constant HD_DATA_TYPE : string := BINARY;
constant DENSE : string := 0;
constant SPARSE : string := 1;
constant HD_MODE : string := DENSE;
constant SIMI_COS : string := 0;
constant SIMI_DPROD : string := 1;
constant SIMI_HAM : string := 2;
constant HD_SIMI_METHOD : string := SIMI_HAM;
constant APPROX_SQRT_ON_HW : string := 0;
constant APPROX_SQRT_ON_MODEL : string := 0;
constant HD_SIMI_W_BITS : string := 32;
constant LINEAR : string := 0;
constant APPROX : string := 1;
constant THERMOMETER : string := 2;
constant HD_LV_TYPE : string := APPROX;
constant HD_LV_LEN : string := 21;
constant SPARSITY_FACTOR_X10 : string := 5;
constant PROBLEM_TYPE_CLASSIFICATION : string := 0;
constant PROBLEM_TYPE_CLUSTERING : string := 1;
constant PROBLEM_TYPE_REGRESSION : string := 2;
constant PROBLEM_TYPE : string := PROBLEM_TYPE_CLASSIFICATION;
constant DI_M_STREAM : string := 0;
constant DI_M_PARTIAL_PARALLEL : string := 1;
constant DI_M_PARALLEL : string := 2;
constant IN_DATA_MODE : string := DI_M_STREAM;
constant AXI_CNTR_PORT_EN : string := 0;
constant PARALLELISM_FEATURES : string := 1;
constant PARALLELISM_CLASS : string := 1;
constant DI_PARALLEL_W_BITS : string := 64;
constant FRAME_SIZE_MIN : string := 64;
constant DI_QUANT_BITS : string := 6;
constant HD_DATA_W_BITS : string := 1;
constant BV_M_INT_MEM : string := 0;
constant BV_M_EXT : string := 1;
constant BV_M_PERMUTATION : string := 2;
constant BV_M_RND_GEN : string := 3;
constant BV_MODE : string := BV_M_INT_MEM;
constant BV_DATA_W_BITS : string := 1;
constant BV_IN_DATA_W_BITS : string := 64;
constant BV_RND_GEN_W_BITS : string := 64;
constant LV_M_INT_MEM : string := 0;
constant LV_M_EXT : string := 1;
constant LV_M_LOGIC : string := 2;
constant LV_M_HDL_GEN : string := 3;
constant LV_MODE : string := LV_M_INT_MEM;
constant LV_DATA_W_BITS : string := 1;
constant LV_IN_DATA_W_BITS : string := 64;
constant LV_M_APPROX_RND_GEN_W_BITS : string := 64;
constant CV_M_INT_MEM : string := 0;
constant CV_M_EXT : string := 1;
constant CV_M_HDL_GEN : string := 2;
constant CV_MODE : string := CV_M_INT_MEM;
constant CV_DATA_W_BITS : string := 1;
constant CV_IN_DATA_W_BITS : string := 64;
constant DI_FEATUREID_W_BITS : string := 10;
constant DI_FRAMEID_W_BITS : string := 10;
constant DO_CLASS_W_BITS : string := 6;
constant DO_STATUS_W_BITS : string := 5;
constant HD_BUNDLE_W_BITS : string := 32;
constant ENCODING_RECORD : string := 0;
constant ENCODING_NGRAM : string := 1;
constant ENCODING_TECHNIQUE : string := ENCODING_RECORD;
constant N_GRAM_SIZE : string := 4;
constant N_GRAM : string := 1;
constant CLIPPING_DISABLE : string := 0;
constant CLIPPING_BINARY : string := 1;
constant CLIPPING_TERNARY : string := 2;
constant CLIPPING_QUANTIZED : string := 3;
constant CLIPPING_POWERTWO : string := 4;
constant CLIPPING_QUANTIZED_POWERTWO : string := 5;
constant CLIPPING_THRESHOLD : string := 6;
constant CLIPPING_ENCODING : string := CLIPPING_BINARY;
constant CLIPPING_CLASS : string := CLIPPING_BINARY;
constant CLIPPING_BINARY_FOR_VALUE_EQ_HALF_HD_DIM_USE_TOGGLING : string := 0;
constant CLIPPING_BINARY_FOR_VALUE_EQ_HALF_HD_DIM_SET_ZERO : string := 1;
constant CLIPPING_BINARY_METHOD_FOR_VALUE_EQ_HALF_HD_DIM : string := CLIPPING_BINARY_FOR_VALUE_EQ_HALF_HD_DIM_SET_ZERO;
constant HW_CLIPPING_AFTER_TRAIN : string := 0;
constant QUANT_MIN : string := 0;
constant QUANT_MAX : string := 1024;
constant LR_CONSTANT : string := 0;
constant LR_ITER : string := 1;
constant LR_DATA : string := 2;
constant LR_HYBRID : string := 3;
constant LR_DECAY : string := LR_CONSTANT;
constant MAX_LEARNING_RATE : string := 50;
constant BETA_LR : string := 3;
constant RETRAIN : string := 0;
constant VITIS_HLS_XILINX_PATH : string := "C:/Xilinx/Vitis_HLS/2023.1/bin/vitis_hls.bat";
constant VIVADO_XILINX_PATH : string := "C:/Xilinx/Vivado/2023.1/bin/vivado.bat";
constant VITIS_XILINX_PATH : string := "C:/Xilinx/Vitis/2023.1/bin/vitis.bat";
