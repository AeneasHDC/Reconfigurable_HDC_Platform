----
 -- @file level_hvec_gen_hdl.hpp
 -- @brief This script generates HDL code for generating high-dimensional LEVEL vectors.
 -- It is a novel method; for more information, please refer to our paper.
 --
 -- @author Saeid Jamili and Marco Angioli
 -- @note Author names are listed in alphabetical order.
 -- @email <saeid.jamili@uniroma1.it>
 -- @email <marco.angioli@uniroma1.it>
 --
 -- @contributors
 --
 -- @date Created: 24th July 2023
 -- @date Last Updated: 23th August 2023
 --
 -- @version 1.0.0
 --
 -- @institute Sapienza University of Rome
 -- @cite https://doi.org/10.xxxx/yyyyy
 --
 -- @section DEPENDENCIES
 -- - Dependency1: Description or version details.
 -- - Dependency2: Description or version details.
 --
 -- @section LICENSE
 -- This file is part of the Aeneas HyperCompute Platform.
 --
 -- Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 --
 -- @section CHANGELOG
 -- @version 1.0.0-dev - 23th August 2023
 -- - Initial release
 --
 -- @todo
 -- - Complete level vector generator function
 -- - Add training
 --
 -- @see
 -- -
 -- -
 -- -
 --
 --

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity level_vec_gen is
    Port ( level_vec_out : out  STD_LOGIC_VECTOR (63 downto 0);
           frame_index : in  STD_LOGIC_VECTOR (2 downto 0);
           frame_id : in  STD_LOGIC_VECTOR (4 downto 0));
end level_vec_gen;

architecture Behavioral of level_vec_gen is
begin
    process (frame_index, frame_id)
    begin
        -- Update this function to match your requirements
        case frame_index is
            when "000" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0110101000011000111110101101110110100100010101110101000000111111";
                    when "00001" => level_vec_out <= "0110101000011000111110101101110110100100010101110101000000111111";
                    when "00010" => level_vec_out <= "0110111000011000111110101101110110100100010101110101100001111111";
                    when "00011" => level_vec_out <= "0110111101011000111110101101110110100100010101110101100001111111";
                    when "00100" => level_vec_out <= "0110111101011000111110101101110110100100010101110101100001111111";
                    when "00101" => level_vec_out <= "1110111101011000111110101101110110100100010101110101100001111111";
                    when "00110" => level_vec_out <= "1110111101011000111110101101110110100100010101110101100001111111";
                    when "00111" => level_vec_out <= "1110111111011000111111101101110110101100010101110101100001111111";
                    when "01000" => level_vec_out <= "1110111111011000111111101101110110101100010101110101100001111111";
                    when "01001" => level_vec_out <= "1110111111011000111111101101110110101100010101110101101001111111";
                    when "01010" => level_vec_out <= "1110111111011000111111101101110110101100010101110101101001111111";
                    when "01011" => level_vec_out <= "1110111111011010111111101101110110101100011101110101101001111111";
                    when "01100" => level_vec_out <= "1110111111011010111111101101110110101100011101111101101001111111";
                    when "01101" => level_vec_out <= "1110111111011010111111101101110110101100011101111101111001111111";
                    when "01110" => level_vec_out <= "1110111111011010111111101101110110101100011101111101111001111111";
                    when "01111" => level_vec_out <= "1110111111011110111111101101110110101100011111111101111001111111";
                    when "10000" => level_vec_out <= "1110111111011110111111111101110110101100011111111101111001111111";
                    when "10001" => level_vec_out <= "1111111111011110111111111101110110101100011111111101111001111111";
                    when "10010" => level_vec_out <= "1111111111011110111111111101110110101100011111111111111001111111";
                    when "10011" => level_vec_out <= "1111111111011110111111111101110110101100011111111111111001111111";
                    when "10100" => level_vec_out <= "1111111111011110111111111101110110101110011111111111111001111111";
                    when "10101" => level_vec_out <= "1111111111011110111111111101110110101110011111111111111001111111";
                    when "10110" => level_vec_out <= "1111111111011110111111111101110111101110011111111111111001111111";
                    when "10111" => level_vec_out <= "1111111111011110111111111101110111101111011111111111111001111111";
                    when "11000" => level_vec_out <= "1111111111011110111111111101110111101111011111111111111001111111";
                    when "11001" => level_vec_out <= "1111111111111110111111111101110111101111011111111111111001111111";
                    when "11010" => level_vec_out <= "1111111111111110111111111101110111101111011111111111111101111111";
                    when "11011" => level_vec_out <= "1111111111111110111111111101110111101111011111111111111101111111";
                    when "11100" => level_vec_out <= "1111111111111111111111111101110111101111011111111111111101111111";
                    when "11101" => level_vec_out <= "1111111111111111111111111111111111101111011111111111111101111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111101111011111111111111101111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111101111011111111111111101111111";
                when others => null;
                end case;
            when "001" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0011110001000100101010000000010110101101010110011100110001101111";
                    when "00001" => level_vec_out <= "0011110001001101101010010001010110101101010110011100110011101111";
                    when "00010" => level_vec_out <= "0011110001001101101010010001010110101101110110011100110011101111";
                    when "00011" => level_vec_out <= "0111110001001101101010010001010110101101110110011100110011101111";
                    when "00100" => level_vec_out <= "0111110001001101101010010001010110101101110110011100110011101111";
                    when "00101" => level_vec_out <= "0111110001001101101010010001110110101101110110011100110011101111";
                    when "00110" => level_vec_out <= "0111110001001101101010110101110110101101110110011100110011101111";
                    when "00111" => level_vec_out <= "0111110001001111101010110101110110101101111110011100110011101111";
                    when "01000" => level_vec_out <= "0111110001001111101110110101110110101101111110011100110111101111";
                    when "01001" => level_vec_out <= "0111110001001111101110110101110110101111111110011100110111101111";
                    when "01010" => level_vec_out <= "0111110011001111101110110101110110101111111110011100110111101111";
                    when "01011" => level_vec_out <= "0111110011001111101110110101110111101111111110011100110111101111";
                    when "01100" => level_vec_out <= "0111110011001111101110110101110111101111111110011100110111101111";
                    when "01101" => level_vec_out <= "0111110011001111101110110101111111101111111110111100110111101111";
                    when "01110" => level_vec_out <= "0111110011001111101110110101111111101111111110111100110111101111";
                    when "01111" => level_vec_out <= "0111110011001111111110110101111111101111111110111100111111101111";
                    when "10000" => level_vec_out <= "0111110011001111111110110101111111101111111110111100111111101111";
                    when "10001" => level_vec_out <= "0111111011011111111110110101111111101111111110111100111111101111";
                    when "10010" => level_vec_out <= "0111111011011111111110110101111111101111111110111101111111101111";
                    when "10011" => level_vec_out <= "0111111011011111111110110101111111101111111110111101111111111111";
                    when "10100" => level_vec_out <= "0111111011011111111110110101111111101111111110111101111111111111";
                    when "10101" => level_vec_out <= "0111111011011111111111110111111111101111111110111101111111111111";
                    when "10110" => level_vec_out <= "0111111011011111111111110111111111101111111110111101111111111111";
                    when "10111" => level_vec_out <= "1111111011011111111111110111111111101111111110111101111111111111";
                    when "11000" => level_vec_out <= "1111111011011111111111110111111111111111111110111101111111111111";
                    when "11001" => level_vec_out <= "1111111011011111111111110111111111111111111110111101111111111111";
                    when "11010" => level_vec_out <= "1111111011011111111111110111111111111111111111111101111111111111";
                    when "11011" => level_vec_out <= "1111111011011111111111110111111111111111111111111101111111111111";
                    when "11100" => level_vec_out <= "1111111011011111111111110111111111111111111111111101111111111111";
                    when "11101" => level_vec_out <= "1111111011011111111111110111111111111111111111111111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "010" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1001010000000001011000110001100001100100000011111111101101000011";
                    when "00001" => level_vec_out <= "1001010000000001011000110001110001100100000011111111101101000011";
                    when "00010" => level_vec_out <= "1001010000000001011000110001110001100100000011111111101101000011";
                    when "00011" => level_vec_out <= "1001010000000001011000110011110001100101000011111111101101000011";
                    when "00100" => level_vec_out <= "1101010000000001011000110011110001100101000011111111101101000011";
                    when "00101" => level_vec_out <= "1101010000000001011000110111110001100101000011111111101101001011";
                    when "00110" => level_vec_out <= "1101010010000001011000110111110001100101000011111111101101001011";
                    when "00111" => level_vec_out <= "1101010010000001011000110111110001100101000011111111101101001011";
                    when "01000" => level_vec_out <= "1101010010000001011000110111110001100101000011111111101101001011";
                    when "01001" => level_vec_out <= "1101010010010001011000110111110001100101000011111111101101001011";
                    when "01010" => level_vec_out <= "1101010010010001011010110111110001100101000011111111101101001011";
                    when "01011" => level_vec_out <= "1101010010110001011010110111110001100101000011111111101101001011";
                    when "01100" => level_vec_out <= "1101010010110001011010110111110001100111000011111111101101001011";
                    when "01101" => level_vec_out <= "1101010010110001011010110111110001100111000011111111101101001011";
                    when "01110" => level_vec_out <= "1101010010110101011010110111110001100111000011111111101101011011";
                    when "01111" => level_vec_out <= "1101010010110101011010110111110001100111000011111111101101011011";
                    when "10000" => level_vec_out <= "1101010010110101011010110111110001101111000011111111101101011011";
                    when "10001" => level_vec_out <= "1101010010110101011010110111110001101111000011111111111101011011";
                    when "10010" => level_vec_out <= "1101010010110101011010110111110001101111000111111111111101111011";
                    when "10011" => level_vec_out <= "1101010010110101011010110111110001101111000111111111111101111111";
                    when "10100" => level_vec_out <= "1101011010110101011010110111110001111111010111111111111101111111";
                    when "10101" => level_vec_out <= "1111011010110101011010110111111001111111010111111111111101111111";
                    when "10110" => level_vec_out <= "1111011010110101011010110111111001111111010111111111111101111111";
                    when "10111" => level_vec_out <= "1111011010110101011010110111111001111111010111111111111101111111";
                    when "11000" => level_vec_out <= "1111011010110101011011110111111001111111010111111111111111111111";
                    when "11001" => level_vec_out <= "1111111110110101011011110111111001111111010111111111111111111111";
                    when "11010" => level_vec_out <= "1111111110110101011011110111111001111111010111111111111111111111";
                    when "11011" => level_vec_out <= "1111111110110101011111110111111001111111110111111111111111111111";
                    when "11100" => level_vec_out <= "1111111110110101011111110111111101111111110111111111111111111111";
                    when "11101" => level_vec_out <= "1111111110110101011111110111111101111111110111111111111111111111";
                    when "11110" => level_vec_out <= "1111111110110101011111110111111101111111110111111111111111111111";
                    when "11111" => level_vec_out <= "1111111110111101111111110111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "011" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0111000001100010100101001001100001011111000111100100010100010111";
                    when "00001" => level_vec_out <= "0111000001100010100101001001101001011111000111100100010100010111";
                    when "00010" => level_vec_out <= "0111000011100010100101001001101001011111000111100100010100010111";
                    when "00011" => level_vec_out <= "0111000011100010100101001001101001011111000111100100010100010111";
                    when "00100" => level_vec_out <= "0111000011100010100101001101101001011111010111100100010100010111";
                    when "00101" => level_vec_out <= "0111000011100010100101001101101001011111010111100100010100010111";
                    when "00110" => level_vec_out <= "0111000111100010100101001101101001011111010111100100010100010111";
                    when "00111" => level_vec_out <= "0111000111100010100101001101101001011111010111100100010100010111";
                    when "01000" => level_vec_out <= "0111000111100010100101001101101001011111011111110100010100010111";
                    when "01001" => level_vec_out <= "0111000111100010110101001111101001011111011111110100010100010111";
                    when "01010" => level_vec_out <= "0111000111100010110111001111101001011111011111110100010100010111";
                    when "01011" => level_vec_out <= "0111000111100011110111001111101001011111011111110100010100011111";
                    when "01100" => level_vec_out <= "0111000111100011110111001111101001011111011111110100010100011111";
                    when "01101" => level_vec_out <= "0111000111100011110111001111101001011111011111110100010110011111";
                    when "01110" => level_vec_out <= "0111000111100011110111001111101011011111111111110100010110011111";
                    when "01111" => level_vec_out <= "0111001111100011110111001111101011011111111111110100010110011111";
                    when "10000" => level_vec_out <= "1111101111100011110111001111101011011111111111110100010110011111";
                    when "10001" => level_vec_out <= "1111101111100011110111001111101011011111111111110100010110011111";
                    when "10010" => level_vec_out <= "1111101111100011110111101111101011011111111111110100010110011111";
                    when "10011" => level_vec_out <= "1111101111100011110111101111101011011111111111110100010110011111";
                    when "10100" => level_vec_out <= "1111101111100011110111101111101011011111111111110100010110011111";
                    when "10101" => level_vec_out <= "1111111111100011110111111111101011111111111111110100010110011111";
                    when "10110" => level_vec_out <= "1111111111100011110111111111101011111111111111110100011110011111";
                    when "10111" => level_vec_out <= "1111111111110011110111111111101011111111111111110100011110011111";
                    when "11000" => level_vec_out <= "1111111111110011111111111111101011111111111111110101011110011111";
                    when "11001" => level_vec_out <= "1111111111111011111111111111111011111111111111110101011111011111";
                    when "11010" => level_vec_out <= "1111111111111011111111111111111011111111111111110101011111011111";
                    when "11011" => level_vec_out <= "1111111111111011111111111111111011111111111111111101011111011111";
                    when "11100" => level_vec_out <= "1111111111111011111111111111111011111111111111111101011111011111";
                    when "11101" => level_vec_out <= "1111111111111011111111111111111111111111111111111101011111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111111111111101011111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "100" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0001101100011100001101111011010110001001001000010101111011101100";
                    when "00001" => level_vec_out <= "0001101100011100001101111011010110001001001000010101111011101100";
                    when "00010" => level_vec_out <= "0001101100011100001101111011010110001001001000010101111011101100";
                    when "00011" => level_vec_out <= "0001111100011100001101111011011110001001001000010101111011101100";
                    when "00100" => level_vec_out <= "0001111100011100001101111011111110001001001000010101111011101101";
                    when "00101" => level_vec_out <= "0001111100011100001101111011111110001001001000010101111011101101";
                    when "00110" => level_vec_out <= "0001111100011101001101111011111110001001001010010101111011101101";
                    when "00111" => level_vec_out <= "0001111100011101001101111011111110001001011010010101111111101101";
                    when "01000" => level_vec_out <= "0001111100011101001101111011111110001001011010011101111111101101";
                    when "01001" => level_vec_out <= "0111111100011101001101111011111110001001011010011101111111101101";
                    when "01010" => level_vec_out <= "0111111100011101001101111011111110101001011010011101111111111101";
                    when "01011" => level_vec_out <= "0111111100011101001101111011111110101001011010011101111111111101";
                    when "01100" => level_vec_out <= "0111111100011111101101111111111110101001011010011101111111111101";
                    when "01101" => level_vec_out <= "0111111110011111101111111111111110101001111010011101111111111101";
                    when "01110" => level_vec_out <= "0111111110011111101111111111111110101001111010011111111111111101";
                    when "01111" => level_vec_out <= "0111111110011111101111111111111110101001111010011111111111111101";
                    when "10000" => level_vec_out <= "0111111110011111101111111111111110101001111010011111111111111101";
                    when "10001" => level_vec_out <= "0111111110011111101111111111111110101001111110011111111111111101";
                    when "10010" => level_vec_out <= "0111111110011111101111111111111110101001111110011111111111111101";
                    when "10011" => level_vec_out <= "0111111110011111111111111111111110101001111110011111111111111101";
                    when "10100" => level_vec_out <= "0111111110011111111111111111111110101101111110011111111111111101";
                    when "10101" => level_vec_out <= "0111111110011111111111111111111110101101111110011111111111111101";
                    when "10110" => level_vec_out <= "0111111110011111111111111111111111101101111110011111111111111101";
                    when "10111" => level_vec_out <= "0111111110011111111111111111111111101101111110011111111111111101";
                    when "11000" => level_vec_out <= "0111111110011111111111111111111111111101111110011111111111111111";
                    when "11001" => level_vec_out <= "0111111110011111111111111111111111111101111110011111111111111111";
                    when "11010" => level_vec_out <= "0111111110011111111111111111111111111101111110111111111111111111";
                    when "11011" => level_vec_out <= "0111111110011111111111111111111111111111111110111111111111111111";
                    when "11100" => level_vec_out <= "1111111111011111111111111111111111111111111110111111111111111111";
                    when "11101" => level_vec_out <= "1111111111011111111111111111111111111111111110111111111111111111";
                    when "11110" => level_vec_out <= "1111111111011111111111111111111111111111111110111111111111111111";
                    when "11111" => level_vec_out <= "1111111111011111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "101" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0000011001001000001010011110010111101111101000100010100110010111";
                    when "00001" => level_vec_out <= "0000011001001000001010011110010111101111101000100010110110010111";
                    when "00010" => level_vec_out <= "0000011001001000001010011110010111101111101000100010110110010111";
                    when "00011" => level_vec_out <= "0000011001001000001010011110010111101111101000100110110110010111";
                    when "00100" => level_vec_out <= "0000011001001000001010011110010111101111101000100111110110010111";
                    when "00101" => level_vec_out <= "0000111001001000001010011110010111101111101000100111110110010111";
                    when "00110" => level_vec_out <= "0000111001001000001010011110010111101111101000100111110110010111";
                    when "00111" => level_vec_out <= "0000111001001000101010011110010111101111101000100111110110010111";
                    when "01000" => level_vec_out <= "0000111001001000101010011110010111101111101000100111110111011111";
                    when "01001" => level_vec_out <= "0000111001001000101010011110010111101111101000100111110111011111";
                    when "01010" => level_vec_out <= "0000111001001100101010011110010111101111101000100111110111011111";
                    when "01011" => level_vec_out <= "0000111001001100101010011110010111101111101001100111110111011111";
                    when "01100" => level_vec_out <= "0001111001001100101010011110011111101111101001100111110111011111";
                    when "01101" => level_vec_out <= "0001111001001100101010011110011111101111101001100111110111011111";
                    when "01110" => level_vec_out <= "0001111001001100101010011110011111101111101101100111110111011111";
                    when "01111" => level_vec_out <= "0001111101001100101010011110111111101111101101110111110111011111";
                    when "10000" => level_vec_out <= "0001111101011100101010011110111111101111101111110111110111011111";
                    when "10001" => level_vec_out <= "0001111101011100111011011110111111101111101111110111110111011111";
                    when "10010" => level_vec_out <= "0001111111011100111011011110111111101111101111110111110111011111";
                    when "10011" => level_vec_out <= "0101111111011101111011011110111111101111101111110111110111011111";
                    when "10100" => level_vec_out <= "0111111111011101111011011110111111101111101111110111110111011111";
                    when "10101" => level_vec_out <= "0111111111011101111011011110111111101111101111110111110111011111";
                    when "10110" => level_vec_out <= "0111111111111111111011011110111111101111101111110111111111011111";
                    when "10111" => level_vec_out <= "0111111111111111111011011110111111101111111111110111111111011111";
                    when "11000" => level_vec_out <= "0111111111111111111011011110111111101111111111110111111111011111";
                    when "11001" => level_vec_out <= "0111111111111111111011011110111111101111111111110111111111011111";
                    when "11010" => level_vec_out <= "1111111111111111111011111110111111101111111111110111111111011111";
                    when "11011" => level_vec_out <= "1111111111111111111011111110111111101111111111110111111111011111";
                    when "11100" => level_vec_out <= "1111111111111111111011111111111111111111111111110111111111011111";
                    when "11101" => level_vec_out <= "1111111111111111111011111111111111111111111111111111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111011111111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111011111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "110" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1111011111001010001111011111010000011111111001101100011111011000";
                    when "00001" => level_vec_out <= "1111011111001010001111011111010000011111111001101100011111011000";
                    when "00010" => level_vec_out <= "1111011111001011001111011111010000011111111001101100011111011101";
                    when "00011" => level_vec_out <= "1111011111001011001111011111010000011111111001101100011111011101";
                    when "00100" => level_vec_out <= "1111011111001011001111011111010000011111111001101100011111011101";
                    when "00101" => level_vec_out <= "1111011111001111001111011111010000011111111001101100011111011101";
                    when "00110" => level_vec_out <= "1111011111001111001111011111010100011111111001111100011111011101";
                    when "00111" => level_vec_out <= "1111011111001111001111011111010100011111111001111100011111011101";
                    when "01000" => level_vec_out <= "1111011111001111001111011111010100011111111001111100111111011101";
                    when "01001" => level_vec_out <= "1111011111001111001111011111010100011111111001111110111111011101";
                    when "01010" => level_vec_out <= "1111011111001111001111011111010100011111111001111110111111011101";
                    when "01011" => level_vec_out <= "1111011111001111101111011111010100011111111001111110111111011101";
                    when "01100" => level_vec_out <= "1111011111001111101111011111010100011111111001111110111111011101";
                    when "01101" => level_vec_out <= "1111011111001111101111011111010100011111111001111110111111011101";
                    when "01110" => level_vec_out <= "1111011111001111101111011111010100011111111001111110111111011101";
                    when "01111" => level_vec_out <= "1111011111001111101111011111010100011111111001111110111111011101";
                    when "10000" => level_vec_out <= "1111011111011111101111011111010100011111111001111110111111011101";
                    when "10001" => level_vec_out <= "1111011111011111101111011111010100011111111001111110111111011101";
                    when "10010" => level_vec_out <= "1111011111011111101111011111010100111111111001111110111111011101";
                    when "10011" => level_vec_out <= "1111011111011111101111011111010100111111111011111110111111011111";
                    when "10100" => level_vec_out <= "1111011111011111101111011111010100111111111011111110111111011111";
                    when "10101" => level_vec_out <= "1111011111011111101111011111010100111111111011111111111111011111";
                    when "10110" => level_vec_out <= "1111111111011111101111011111010100111111111011111111111111011111";
                    when "10111" => level_vec_out <= "1111111111011111101111011111110100111111111011111111111111011111";
                    when "11000" => level_vec_out <= "1111111111011111101111011111110100111111111011111111111111011111";
                    when "11001" => level_vec_out <= "1111111111011111101111011111110100111111111011111111111111011111";
                    when "11010" => level_vec_out <= "1111111111111111101111011111110101111111111011111111111111011111";
                    when "11011" => level_vec_out <= "1111111111111111111111011111110101111111111111111111111111011111";
                    when "11100" => level_vec_out <= "1111111111111111111111111111110101111111111111111111111111011111";
                    when "11101" => level_vec_out <= "1111111111111111111111111111110101111111111111111111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111110111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "111" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1111011010111000110110000010101010011111001110001011001000111010";
                    when "00001" => level_vec_out <= "1111011010111000110110000010101010011111001110001011001000111010";
                    when "00010" => level_vec_out <= "1111011010111000110110000010101010011111001110001011001000111010";
                    when "00011" => level_vec_out <= "1111011010111000110110000010101010011111001110001011001000111010";
                    when "00100" => level_vec_out <= "1111011010111000110110000110101010011111001110001011001001111010";
                    when "00101" => level_vec_out <= "1111011010111000110110000110101110011111001110101011001001111010";
                    when "00110" => level_vec_out <= "1111011010111000110110000110101110011111001110101011001001111010";
                    when "00111" => level_vec_out <= "1111011010111000110110000110101110011111001110101011001001111010";
                    when "01000" => level_vec_out <= "1111011010111000110110000110101110011111001110101011001001111010";
                    when "01001" => level_vec_out <= "1111011010111000110110000110101110011111001110101011001001111010";
                    when "01010" => level_vec_out <= "1111011010111000110110010110101110011111001111101011001001111010";
                    when "01011" => level_vec_out <= "1111011010111000110110010110101110011111001111101011001001111010";
                    when "01100" => level_vec_out <= "1111011010111000110110010110101110011111001111101011001001111110";
                    when "01101" => level_vec_out <= "1111011010111000110110010110101110011111001111101011011001111110";
                    when "01110" => level_vec_out <= "1111011010111000110111010110101110011111001111111011011001111110";
                    when "01111" => level_vec_out <= "1111011010111000110111010110101110011111001111111011011001111110";
                    when "10000" => level_vec_out <= "1111011010111000110111010110101110111111001111111011011001111110";
                    when "10001" => level_vec_out <= "1111011110111000110111010110101110111111001111111011011001111110";
                    when "10010" => level_vec_out <= "1111011110111000110111010110101110111111001111111111011001111110";
                    when "10011" => level_vec_out <= "1111011110111000110111010110101110111111101111111111011001111110";
                    when "10100" => level_vec_out <= "1111011110111100110111011110101110111111101111111111011001111110";
                    when "10101" => level_vec_out <= "1111011110111100110111011110101110111111101111111111011001111110";
                    when "10110" => level_vec_out <= "1111011110111100110111011110101111111111101111111111011001111110";
                    when "10111" => level_vec_out <= "1111011110111111110111111110101111111111101111111111011001111110";
                    when "11000" => level_vec_out <= "1111011110111111110111111110101111111111101111111111011001111111";
                    when "11001" => level_vec_out <= "1111011111111111110111111110101111111111101111111111011101111111";
                    when "11010" => level_vec_out <= "1111011111111111111111111110101111111111101111111111011101111111";
                    when "11011" => level_vec_out <= "1111111111111111111111111110101111111111111111111111011101111111";
                    when "11100" => level_vec_out <= "1111111111111111111111111110111111111111111111111111011101111111";
                    when "11101" => level_vec_out <= "1111111111111111111111111110111111111111111111111111011101111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when others => null;
        end case;
    end process;
end Behavioral;