/**
 * @file level_hvec_gen_hdl.hpp
 * @brief This script generates HDL code for generating high-dimensional LEVEL vectors.
 * It is a novel method; for more information, please refer to our paper.
 *
 * @author Saeid Jamili and Marco Angioli
 * @note Author names are listed in alphabetical order.
 * @email <saeid.jamili@uniroma1.it>
 * @email <marco.angioli@uniroma1.it>
 *
 * @contributors
 *
 * @date Created: 24th July 2023
 * @date Last Updated: 23th August 2023
 *
 * @version 1.0.0
 *
 * @institute Sapienza University of Rome
 * @cite https://doi.org/10.xxxx/yyyyy
 *
 * @section DEPENDENCIES
 * - Dependency1: Description or version details.
 * - Dependency2: Description or version details.
 *
 * @section LICENSE
 * This file is part of the Aeneas HyperCompute Platform.
 *
 * Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 *
 * @section CHANGELOG
 * @version 1.0.0-dev - 23th August 2023
 * - Initial release
 *
 * @todo
 * - Complete level vector generator function
 * - Add training
 *
 * @see
 * -
 * -
 * -
 *
 */

module level_vec_gen (
    output reg [63:0] level_vec_out,
    input [2:0] frame_index,
    input [4:0] frame_id
);
    always @(*) begin
        // Update this function to match your requirements
        case (frame_index)
            0: begin
                case (frame_id)
                    0: level_vec_out = 64'b1000100110001011101101101111001110000110111001011001010000010000;
                    1: level_vec_out = 64'b1000100110001011101101101111001110000110111001011001010000010001;
                    2: level_vec_out = 64'b1000100110001011101101101111001110000110111001011001010000010001;
                    3: level_vec_out = 64'b1000100111001011101111101111011111000110111001011001010000010011;
                    4: level_vec_out = 64'b1000100111001011101111101111011111000110111001011001010000010011;
                    5: level_vec_out = 64'b1000100111001011101111101111011111000110111101011001010000010011;
                    6: level_vec_out = 64'b1000100111001011101111111111011111000110111101011001010000010011;
                    7: level_vec_out = 64'b1010100111001011101111111111011111000110111101011001010000010011;
                    8: level_vec_out = 64'b1010100111001011101111111111011111000111111101011001010000010011;
                    9: level_vec_out = 64'b1011100111001011101111111111011111000111111101011001010000010011;
                    10: level_vec_out = 64'b1011100111001011101111111111011111000111111101011001010000011011;
                    11: level_vec_out = 64'b1011100111001011101111111111011111000111111101011001010000011011;
                    12: level_vec_out = 64'b1011100111001011101111111111011111000111111101011001010100011011;
                    13: level_vec_out = 64'b1011100111001011101111111111011111000111111101011001010100111011;
                    14: level_vec_out = 64'b1011100111001011101111111111011111000111111101111001010100111111;
                    15: level_vec_out = 64'b1011100111001011101111111111011111010111111101111001010110111111;
                    16: level_vec_out = 64'b1011100111001011101111111111011111010111111101111001010110111111;
                    17: level_vec_out = 64'b1011100111001011101111111111011111010111111101111001010111111111;
                    18: level_vec_out = 64'b1011100111001011101111111111011111010111111101111001110111111111;
                    19: level_vec_out = 64'b1011100111001011101111111111011111011111111111111011110111111111;
                    20: level_vec_out = 64'b1011100111001011101111111111011111011111111111111011110111111111;
                    21: level_vec_out = 64'b1011100111001011111111111111011111011111111111111011110111111111;
                    22: level_vec_out = 64'b1011100111001011111111111111011111011111111111111011110111111111;
                    23: level_vec_out = 64'b1011100111001011111111111111011111011111111111111011111111111111;
                    24: level_vec_out = 64'b1111100111001011111111111111011111011111111111111011111111111111;
                    25: level_vec_out = 64'b1111100111001011111111111111011111111111111111111011111111111111;
                    26: level_vec_out = 64'b1111100111001011111111111111011111111111111111111011111111111111;
                    27: level_vec_out = 64'b1111100111001011111111111111011111111111111111111011111111111111;
                    28: level_vec_out = 64'b1111100111101111111111111111011111111111111111111011111111111111;
                    29: level_vec_out = 64'b1111100111101111111111111111011111111111111111111011111111111111;
                    30: level_vec_out = 64'b1111110111101111111111111111011111111111111111111111111111111111;
                    31: level_vec_out = 64'b1111110111101111111111111111011111111111111111111111111111111111;
                endcase
            end
            1: begin
                case (frame_id)
                    0: level_vec_out = 64'b1001010001110010001111001010001010011001110111111001100100101110;
                    1: level_vec_out = 64'b1001010001110010001111001010001010011101110111111001100100101110;
                    2: level_vec_out = 64'b1011010001110010001111001010001010011101110111111001100110101110;
                    3: level_vec_out = 64'b1011010001110010001111001010001010011101110111111001100110101110;
                    4: level_vec_out = 64'b1111010011110010001111001010001010011101110111111001100110101110;
                    5: level_vec_out = 64'b1111010011110010001111001010001010011101110111111001100110101110;
                    6: level_vec_out = 64'b1111010011110010001111001010001010011101110111111001101110101110;
                    7: level_vec_out = 64'b1111010011110110001111001010001010011101110111111011101110101110;
                    8: level_vec_out = 64'b1111110011110110001111001010001010011101110111111011111110101110;
                    9: level_vec_out = 64'b1111110011110110001111001010001010011101110111111011111110101110;
                    10: level_vec_out = 64'b1111111011111110001111001010001010011101110111111011111110101111;
                    11: level_vec_out = 64'b1111111011111110001111001010001011011101110111111011111110101111;
                    12: level_vec_out = 64'b1111111011111110001111001010001011011101110111111011111110101111;
                    13: level_vec_out = 64'b1111111011111110001111001010001011011101110111111011111110101111;
                    14: level_vec_out = 64'b1111111011111110001111001010001011011101110111111011111110101111;
                    15: level_vec_out = 64'b1111111011111110001111001010001011011101110111111011111110101111;
                    16: level_vec_out = 64'b1111111011111110101111001010101011011101110111111011111110101111;
                    17: level_vec_out = 64'b1111111011111110101111001010101011011101111111111011111110101111;
                    18: level_vec_out = 64'b1111111011111110101111001011101011011101111111111011111110111111;
                    19: level_vec_out = 64'b1111111011111110101111001111101011011101111111111011111110111111;
                    20: level_vec_out = 64'b1111111011111110101111001111101011011101111111111011111110111111;
                    21: level_vec_out = 64'b1111111011111110101111001111101011011101111111111011111111111111;
                    22: level_vec_out = 64'b1111111011111110101111001111101011011101111111111011111111111111;
                    23: level_vec_out = 64'b1111111011111110101111001111101111011101111111111111111111111111;
                    24: level_vec_out = 64'b1111111011111110101111001111101111011101111111111111111111111111;
                    25: level_vec_out = 64'b1111111011111110111111001111101111011101111111111111111111111111;
                    26: level_vec_out = 64'b1111111111111110111111001111101111111101111111111111111111111111;
                    27: level_vec_out = 64'b1111111111111110111111001111101111111101111111111111111111111111;
                    28: level_vec_out = 64'b1111111111111110111111001111101111111111111111111111111111111111;
                    29: level_vec_out = 64'b1111111111111111111111011111101111111111111111111111111111111111;
                    30: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    31: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                endcase
            end
            2: begin
                case (frame_id)
                    0: level_vec_out = 64'b1010010100010001111000110101111101111010011101010111000011100010;
                    1: level_vec_out = 64'b1010010100010001111000110101111101111110011101010111000011100010;
                    2: level_vec_out = 64'b1010010100010001111000110101111101111110011101010111000011100010;
                    3: level_vec_out = 64'b1010010100010001111000110101111101111110011101010111000011100010;
                    4: level_vec_out = 64'b1010010100010001111000110101111101111110011101010111000011100010;
                    5: level_vec_out = 64'b1010110100010001111000110101111101111110011101010111100011100010;
                    6: level_vec_out = 64'b1010110100010001111000110101111101111110011101010111100011100010;
                    7: level_vec_out = 64'b1010110100010001111100110101111101111110011101010111110011100010;
                    8: level_vec_out = 64'b1010110100010001111100110101111101111110011101010111110011100010;
                    9: level_vec_out = 64'b1010110100010001111100111101111101111110011101010111110011100010;
                    10: level_vec_out = 64'b1010110100011001111100111101111101111110011101010111110011100010;
                    11: level_vec_out = 64'b1010110100011001111100111101111101111110011101010111110011100010;
                    12: level_vec_out = 64'b1010110100011001111100111101111101111110011101010111110011100010;
                    13: level_vec_out = 64'b1110110100011011111100111101111101111110011101010111110011100011;
                    14: level_vec_out = 64'b1110111100011011111100111101111101111110011111010111110011100011;
                    15: level_vec_out = 64'b1110111100011011111100111101111101111110011111010111110011100011;
                    16: level_vec_out = 64'b1110111100011011111100111111111101111110011111010111110011100011;
                    17: level_vec_out = 64'b1110111100011011111110111111111101111110011111010111110011100011;
                    18: level_vec_out = 64'b1110111100011011111110111111111101111110011111010111110011100011;
                    19: level_vec_out = 64'b1111111100011011111110111111111101111110011111010111110011100011;
                    20: level_vec_out = 64'b1111111100111011111110111111111101111110011111010111110011100011;
                    21: level_vec_out = 64'b1111111100111011111110111111111101111110011111110111110011110011;
                    22: level_vec_out = 64'b1111111110111011111110111111111101111110011111110111110011111011;
                    23: level_vec_out = 64'b1111111110111011111110111111111101111110011111110111110011111011;
                    24: level_vec_out = 64'b1111111110111011111110111111111101111110011111111111111011111011;
                    25: level_vec_out = 64'b1111111110111011111110111111111101111110011111111111111011111011;
                    26: level_vec_out = 64'b1111111111111011111110111111111111111110011111111111111011111011;
                    27: level_vec_out = 64'b1111111111111011111110111111111111111110111111111111111011111011;
                    28: level_vec_out = 64'b1111111111111011111110111111111111111110111111111111111011111011;
                    29: level_vec_out = 64'b1111111111111011111110111111111111111111111111111111111011111011;
                    30: level_vec_out = 64'b1111111111111111111110111111111111111111111111111111111011111011;
                    31: level_vec_out = 64'b1111111111111111111110111111111111111111111111111111111011111111;
                endcase
            end
            3: begin
                case (frame_id)
                    0: level_vec_out = 64'b0011011101000101101101110010011011000001011111001110111010000110;
                    1: level_vec_out = 64'b0011011101000101101101110010011011100001011111001110111010000111;
                    2: level_vec_out = 64'b0011011101000101101101110010011011100001011111001110111010000111;
                    3: level_vec_out = 64'b0011011101000101101101110010011011100001011111011110111010000111;
                    4: level_vec_out = 64'b0011011101000101101101110010011011100001011111011110111010000111;
                    5: level_vec_out = 64'b0011011101000101101101110010011011101001011111011110111010000111;
                    6: level_vec_out = 64'b0011011101000101101101111010011011101001011111011110111010100111;
                    7: level_vec_out = 64'b0011011101000101111101111010011011101001011111011110111010100111;
                    8: level_vec_out = 64'b0011011101000101111101111010011011101001011111011111111010100111;
                    9: level_vec_out = 64'b0011011101001101111101111010111011101001011111011111111010100111;
                    10: level_vec_out = 64'b0011011101001101111101111010111011101001011111011111111010100111;
                    11: level_vec_out = 64'b0011011101001101111101111010111011101001011111011111111110100111;
                    12: level_vec_out = 64'b0011011101001101111101111010111011101001011111011111111110100111;
                    13: level_vec_out = 64'b0011011101001101111101111010111011101001011111011111111110101111;
                    14: level_vec_out = 64'b0011011101001101111111111010111011101001111111011111111110101111;
                    15: level_vec_out = 64'b1011111101011101111111111010111011101001111111011111111110101111;
                    16: level_vec_out = 64'b1011111101011101111111111010111011101001111111011111111110101111;
                    17: level_vec_out = 64'b1011111101011101111111111010111011101001111111011111111110101111;
                    18: level_vec_out = 64'b1111111101011101111111111011111011101001111111011111111110101111;
                    19: level_vec_out = 64'b1111111101011101111111111011111011101001111111011111111110101111;
                    20: level_vec_out = 64'b1111111101011101111111111011111011101001111111011111111110111111;
                    21: level_vec_out = 64'b1111111101011101111111111011111011101001111111011111111110111111;
                    22: level_vec_out = 64'b1111111101111101111111111011111011101101111111111111111110111111;
                    23: level_vec_out = 64'b1111111101111101111111111011111011101101111111111111111110111111;
                    24: level_vec_out = 64'b1111111101111101111111111011111011101101111111111111111110111111;
                    25: level_vec_out = 64'b1111111101111101111111111111111011101101111111111111111110111111;
                    26: level_vec_out = 64'b1111111101111101111111111111111011101101111111111111111110111111;
                    27: level_vec_out = 64'b1111111101111101111111111111111011101101111111111111111110111111;
                    28: level_vec_out = 64'b1111111101111101111111111111111111101101111111111111111110111111;
                    29: level_vec_out = 64'b1111111111111111111111111111111111101101111111111111111110111111;
                    30: level_vec_out = 64'b1111111111111111111111111111111111101101111111111111111110111111;
                    31: level_vec_out = 64'b1111111111111111111111111111111111111101111111111111111111111111;
                endcase
            end
            4: begin
                case (frame_id)
                    0: level_vec_out = 64'b0100101100101001010010011000001110111110111001000011111000001010;
                    1: level_vec_out = 64'b0100101100101001010010011000001110111110111001100011111000001010;
                    2: level_vec_out = 64'b0101101100101001010010011000001110111110111001100011111000001010;
                    3: level_vec_out = 64'b0101101100101001010010011000001110111110111001100011111000001010;
                    4: level_vec_out = 64'b0101101100101001010010011000001111111110111001100011111000001010;
                    5: level_vec_out = 64'b0101101100101001010010011001001111111110111001100011111000001010;
                    6: level_vec_out = 64'b0101111100101001010110011001001111111110111001100011111000101010;
                    7: level_vec_out = 64'b0101111100101001010110011001001111111110111001100011111000101010;
                    8: level_vec_out = 64'b0101111100101001010110011001001111111110111001100011111000101010;
                    9: level_vec_out = 64'b0101111100101111010110011001001111111110111001100011111000101010;
                    10: level_vec_out = 64'b0101111100101111010110111001001111111110111001100011111000101010;
                    11: level_vec_out = 64'b0101111100101111010110111001001111111110111001100011111000101010;
                    12: level_vec_out = 64'b0101111100101111010110111001001111111111111001100011111000101010;
                    13: level_vec_out = 64'b0101111100101111010110111001001111111111111011100011111000101010;
                    14: level_vec_out = 64'b0101111100101111010110111001001111111111111011100111111000101010;
                    15: level_vec_out = 64'b0101111100101111010110111001001111111111111011100111111000101010;
                    16: level_vec_out = 64'b0101111100101111010110111001001111111111111011110111111000101010;
                    17: level_vec_out = 64'b0101111100101111110110111001001111111111111011111111111001101010;
                    18: level_vec_out = 64'b0101111100101111111110111001001111111111111011111111111001101010;
                    19: level_vec_out = 64'b0101111100101111111110111001001111111111111011111111111001101011;
                    20: level_vec_out = 64'b0101111100101111111110111011101111111111111011111111111001101011;
                    21: level_vec_out = 64'b0101111100101111111110111011101111111111111011111111111001101011;
                    22: level_vec_out = 64'b0101111100101111111110111111101111111111111011111111111011101011;
                    23: level_vec_out = 64'b0101111101101111111111111111101111111111111011111111111011101011;
                    24: level_vec_out = 64'b1101111101101111111111111111101111111111111011111111111011101011;
                    25: level_vec_out = 64'b1101111101101111111111111111101111111111111011111111111011101011;
                    26: level_vec_out = 64'b1111111101101111111111111111101111111111111011111111111011101011;
                    27: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111011101011;
                    28: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111011101011;
                    29: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111011111011;
                    30: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111011;
                    31: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111011;
                endcase
            end
            5: begin
                case (frame_id)
                    0: level_vec_out = 64'b0111110000110100111011111100011110110011100100000110100111010110;
                    1: level_vec_out = 64'b0111110000110100111011111100011110110011100100000110100111010110;
                    2: level_vec_out = 64'b1111110000110100111011111100011110110011100100000110100111010110;
                    3: level_vec_out = 64'b1111110000111100111011111100011110110011100100000110100111010110;
                    4: level_vec_out = 64'b1111110000111100111011111101011110110011100100100110100111010110;
                    5: level_vec_out = 64'b1111110000111100111011111101011110110011100100110110100111010110;
                    6: level_vec_out = 64'b1111110000111101111011111101011110110011100100110110100111010110;
                    7: level_vec_out = 64'b1111110000111101111011111101111110110011100100110110100111010110;
                    8: level_vec_out = 64'b1111111000111101111011111101111110110011100100110110100111010110;
                    9: level_vec_out = 64'b1111111000111101111011111101111110110011100100111110100111010110;
                    10: level_vec_out = 64'b1111111000111101111011111101111110110011100100111110100111010110;
                    11: level_vec_out = 64'b1111111011111101111011111101111110110011100100111110100111010110;
                    12: level_vec_out = 64'b1111111011111101111011111101111110110011100101111110100111010110;
                    13: level_vec_out = 64'b1111111011111101111011111101111110110011100101111110110111010111;
                    14: level_vec_out = 64'b1111111011111101111011111101111110110011100101111110110111010111;
                    15: level_vec_out = 64'b1111111011111101111011111101111110110011101101111110110111010111;
                    16: level_vec_out = 64'b1111111011111101111111111101111110110111101101111110110111010111;
                    17: level_vec_out = 64'b1111111011111101111111111101111110111111101101111110110111010111;
                    18: level_vec_out = 64'b1111111011111101111111111101111110111111101101111110110111010111;
                    19: level_vec_out = 64'b1111111011111101111111111101111110111111101101111110110111110111;
                    20: level_vec_out = 64'b1111111011111101111111111101111110111111101101111111110111110111;
                    21: level_vec_out = 64'b1111111011111101111111111101111110111111111101111111110111110111;
                    22: level_vec_out = 64'b1111111011111101111111111101111110111111111101111111110111110111;
                    23: level_vec_out = 64'b1111111011111101111111111101111110111111111101111111110111110111;
                    24: level_vec_out = 64'b1111111011111101111111111101111110111111111101111111110111110111;
                    25: level_vec_out = 64'b1111111011111101111111111111111110111111111101111111110111110111;
                    26: level_vec_out = 64'b1111111011111101111111111111111110111111111101111111110111111111;
                    27: level_vec_out = 64'b1111111111111101111111111111111110111111111101111111110111111111;
                    28: level_vec_out = 64'b1111111111111101111111111111111110111111111101111111111111111111;
                    29: level_vec_out = 64'b1111111111111101111111111111111110111111111101111111111111111111;
                    30: level_vec_out = 64'b1111111111111101111111111111111111111111111111111111111111111111;
                    31: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                endcase
            end
            6: begin
                case (frame_id)
                    0: level_vec_out = 64'b1111100111011010001001101011010100110111100110101100100010101000;
                    1: level_vec_out = 64'b1111100111011010001001101011010100110111100110101100100010101100;
                    2: level_vec_out = 64'b1111100111011010001001101011010101110111100111101100100010101110;
                    3: level_vec_out = 64'b1111100111011010001001101011010101110111100111101101100010101110;
                    4: level_vec_out = 64'b1111100111011010001001101011110101110111100111101101100010101110;
                    5: level_vec_out = 64'b1111100111011010001001101011110101110111100111101101110110101110;
                    6: level_vec_out = 64'b1111100111011010001001101011110101110111100111101101110110101110;
                    7: level_vec_out = 64'b1111100111011010001001101011110111110111100111101101110110101110;
                    8: level_vec_out = 64'b1111100111011010001001101011110111110111110111111101110110101110;
                    9: level_vec_out = 64'b1111100111011010001001101011110111110111110111111101110110101110;
                    10: level_vec_out = 64'b1111100111011010001001101011110111110111110111111101110110101110;
                    11: level_vec_out = 64'b1111100111011010001001101011110111110111110111111111110110101110;
                    12: level_vec_out = 64'b1111100111111010001101111011110111110111110111111111110110101110;
                    13: level_vec_out = 64'b1111100111111010001101111011110111110111110111111111110110101110;
                    14: level_vec_out = 64'b1111100111111010001101111011110111110111110111111111110110101110;
                    15: level_vec_out = 64'b1111100111111010001101111011110111110111110111111111110110101110;
                    16: level_vec_out = 64'b1111100111111010001111111011110111110111110111111111110110101110;
                    17: level_vec_out = 64'b1111100111111010001111111011110111111111110111111111110110101110;
                    18: level_vec_out = 64'b1111100111111010001111111011110111111111110111111111110110101110;
                    19: level_vec_out = 64'b1111100111111010001111111011110111111111110111111111110110101110;
                    20: level_vec_out = 64'b1111100111111010001111111011110111111111111111111111110110111110;
                    21: level_vec_out = 64'b1111110111111010001111111011110111111111111111111111110110111110;
                    22: level_vec_out = 64'b1111110111111010001111111011110111111111111111111111110110111110;
                    23: level_vec_out = 64'b1111110111111010001111111011110111111111111111111111110110111110;
                    24: level_vec_out = 64'b1111110111111010001111111011110111111111111111111111110110111110;
                    25: level_vec_out = 64'b1111110111111010111111111011110111111111111111111111110111111110;
                    26: level_vec_out = 64'b1111110111111011111111111011110111111111111111111111110111111110;
                    27: level_vec_out = 64'b1111110111111011111111111011110111111111111111111111110111111110;
                    28: level_vec_out = 64'b1111110111111011111111111011110111111111111111111111111111111110;
                    29: level_vec_out = 64'b1111110111111011111111111111111111111111111111111111111111111110;
                    30: level_vec_out = 64'b1111110111111011111111111111111111111111111111111111111111111110;
                    31: level_vec_out = 64'b1111111111111011111111111111111111111111111111111111111111111111;
                endcase
            end
            7: begin
                case (frame_id)
                    0: level_vec_out = 64'b0110000010100110000110101100111000000011100000010101010001010101;
                    1: level_vec_out = 64'b0110000010100110010110101100111000000011100000010101010001010101;
                    2: level_vec_out = 64'b0110000010100110010110101100111000000011100000010101110001010101;
                    3: level_vec_out = 64'b0110000010100110010110101100111000000011100000010101110001010101;
                    4: level_vec_out = 64'b0110100010100110010110101100111000000011100000010101111001010101;
                    5: level_vec_out = 64'b0110100010100110010110101100111000000011100000010101111001010101;
                    6: level_vec_out = 64'b0110100010100110010110101100111000000011100000010101111001010101;
                    7: level_vec_out = 64'b0110100010100110010110101100111000000011100000010101111001010101;
                    8: level_vec_out = 64'b0110110010100110010110101100111000000011100000010101111001010101;
                    9: level_vec_out = 64'b0110110010100110010110101100111010000011100000010101111001010101;
                    10: level_vec_out = 64'b0110110010101110010110101100111010000011100000110101111001010101;
                    11: level_vec_out = 64'b0110110010101110110110101100111010010011100010110101111001010101;
                    12: level_vec_out = 64'b0110110010101111110110101100111010010011100110110101111001010101;
                    13: level_vec_out = 64'b0110110010101111110110101100111010010011100110110101111001010101;
                    14: level_vec_out = 64'b0110110010101111110110101101111010010011100110110101111001010101;
                    15: level_vec_out = 64'b0111110010101111110111101101111010010011100110110101111001010101;
                    16: level_vec_out = 64'b0111110010101111110111101101111010010011100110110101111001011101;
                    17: level_vec_out = 64'b0111110010101111110111101101111010010011100110110101111001011101;
                    18: level_vec_out = 64'b0111110010101111110111111111111010010011100110110101111001011101;
                    19: level_vec_out = 64'b0111110010101111110111111111111010110011100110110101111001011101;
                    20: level_vec_out = 64'b0111111010101111110111111111111010110011100110110101111001011101;
                    21: level_vec_out = 64'b0111111010101111110111111111111010111011100110110101111011011101;
                    22: level_vec_out = 64'b0111111010101111110111111111111110111011100110110101111011011101;
                    23: level_vec_out = 64'b0111111010111111110111111111111110111011101110110101111011111101;
                    24: level_vec_out = 64'b0111111110111111110111111111111110111111101110110111111011111111;
                    25: level_vec_out = 64'b0111111110111111111111111111111110111111101110110111111011111111;
                    26: level_vec_out = 64'b0111111110111111111111111111111110111111111110110111111011111111;
                    27: level_vec_out = 64'b1111111111111111111111111111111110111111111110110111111011111111;
                    28: level_vec_out = 64'b1111111111111111111111111111111110111111111111111111111011111111;
                    29: level_vec_out = 64'b1111111111111111111111111111111110111111111111111111111011111111;
                    30: level_vec_out = 64'b1111111111111111111111111111111110111111111111111111111011111111;
                    31: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                endcase
            end
        endcase
    end
endmodule