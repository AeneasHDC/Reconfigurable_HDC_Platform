// Configuration file for SystemVerilog
`define VERBOS_DISABLE 0;
`define VERBOS_L1 1;
`define VERBOS_L2 2;
`define VERBOS VERBOS_L1;
`define WINDOWS 0;
`define LINUX 1;
`define MAC 2;
`define OS WINDOWS;
`define FPGA 0;
`define MICROCONTROLER 1;
`define SOFT_PROCESSOR 2;
`define DEVICE_TYPE MICROCONTROLER;
`define description "Class Vector Modes and Configurations";
`define TARGET_DEVICE "xczu9eg-ffvb1156-2-e";
`define AMD_ZYBO 0;
`define AMD_ZEDBOARD 1;
`define AMD_ZCU106 2;
`define AMD_ZCU102 3;
`define AMD_VCU108 4;
`define TARGET_BOARD AMD_ZCU102;
`define OP_FREQ 200;
`define USE_VIV_EN 1;
`define VIV_OPT_DEFAULT 0;
`define VIV_OPT_RESOURCE 1;
`define VIV_OPT_SPEED 2;
`define VIV_OPT_PERFORMANCE 3;
`define VIV_OPT_METHOD VIV_OPT_DEFAULT;
`define HLS 0;
`define SYSTEM_VERILOG 1;
`define VHDL 2;
`define VERILOG 3;
`define HDL_LANG HLS;
`define PYTHON 4;
`define MATLAB 5;
`define CPP 6;
`define C 7;
`define RUST 8;
`define MODEL_LANG PYTHON;
`define DS_NAME "CARDIO";
`define DS_SIZE 2126;
`define DS_TRAIN_SIZE 1594;
`define DS_TEST_SIZE 532;
`define DS_VALIDATION_SIZE 500;
`define DS_FEATURE_SIZE 21;
`define DS_DATA_TYPE "FP";
`define DS_DATA_RANGE_MIN 0;
`define DS_DATA_RANGE_MAX 1;
`define DS_CLASSES_SIZE 3;
`define TRAIN_ON_HW 0;
`define RETRAIN_ON_HW 0;
`define EPOCH 1;
`define HD_DIM 512;
`define BINARY 0;
`define BIPOLAR 1;
`define HD_DATA_TYPE BINARY;
`define DENSE 0;
`define SPARSE 1;
`define HD_MODE DENSE;
`define SIMI_COS 0;
`define SIMI_DPROD 1;
`define SIMI_HAM 2;
`define HD_SIMI_METHOD SIMI_HAM;
`define APPROX_SQRT_ON_HW 0;
`define APPROX_SQRT_ON_MODEL 0;
`define HD_SIMI_W_BITS 32;
`define LINEAR 0;
`define APPROX 1;
`define THERMOMETER 2;
`define HD_LV_TYPE LINEAR;
`define HD_LV_LEN 32;
`define SPARSITY_FACTOR_X10 5;
`define PROBLEM_TYPE_CLASSIFICATION 0;
`define PROBLEM_TYPE_CLUSTERING 1;
`define PROBLEM_TYPE_REGRESSION 2;
`define PROBLEM_TYPE PROBLEM_TYPE_CLASSIFICATION;
`define DI_M_STREAM 0;
`define DI_M_PARTIAL_PARALLEL 1;
`define DI_M_PARALLEL 2;
`define IN_DATA_MODE DI_M_STREAM;
`define AXI_CNTR_PORT_EN 0;
`define PARALLELISM_FEATURES 1;
`define PARALLELISM_CLASS 1;
`define DI_PARALLEL_W_BITS 64;
`define FRAME_SIZE_MIN 64;
`define DI_QUANT_BITS 6;
`define HD_DATA_W_BITS 1;
`define BV_M_INT_MEM 0;
`define BV_M_EXT 1;
`define BV_M_PERMUTATION 2;
`define BV_M_RND_GEN 3;
`define BV_MODE BV_M_INT_MEM;
`define BV_DATA_W_BITS 1;
`define BV_IN_DATA_W_BITS 64;
`define BV_RND_GEN_W_BITS 64;
`define LV_M_INT_MEM 0;
`define LV_M_EXT 1;
`define LV_M_LOGIC 2;
`define LV_M_HDL_GEN 3;
`define LV_MODE LV_M_INT_MEM;
`define LV_DATA_W_BITS 1;
`define LV_IN_DATA_W_BITS 64;
`define LV_M_APPROX_RND_GEN_W_BITS 64;
`define CV_M_INT_MEM 0;
`define CV_M_EXT 1;
`define CV_M_HDL_GEN 2;
`define CV_MODE CV_M_INT_MEM;
`define CV_DATA_W_BITS 1;
`define CV_IN_DATA_W_BITS 64;
`define DI_FEATUREID_W_BITS 10;
`define DI_FRAMEID_W_BITS 10;
`define DO_CLASS_W_BITS 6;
`define DO_STATUS_W_BITS 5;
`define HD_BUNDLE_W_BITS 32;
`define ENCODING_RECORD 0;
`define ENCODING_NGRAM 1;
`define ENCODING_TECHNIQUE ENCODING_RECORD;
`define N_GRAM_SIZE 1;
`define N_GRAM 0;
`define CLIPPING_DISABLE 0;
`define CLIPPING_BINARY 1;
`define CLIPPING_TERNARY 2;
`define CLIPPING_QUANTIZED 3;
`define CLIPPING_POWERTWO 4;
`define CLIPPING_QUANTIZED_POWERTWO 5;
`define CLIPPING_THRESHOLD 6;
`define CLIPPING_ENCODING CLIPPING_BINARY;
`define CLIPPING_CLASS CLIPPING_BINARY;
`define CLIPPING_BINARY_FOR_VALUE_EQ_HALF_HD_DIM_USE_TOGGLING 0;
`define CLIPPING_BINARY_FOR_VALUE_EQ_HALF_HD_DIM_SET_ZERO 1;
`define CLIPPING_BINARY_METHOD_FOR_VALUE_EQ_HALF_HD_DIM CLIPPING_BINARY_FOR_VALUE_EQ_HALF_HD_DIM_SET_ZERO;
`define HW_CLIPPING_AFTER_TRAIN 0;
`define QUANT_MIN 0;
`define QUANT_MAX 1;
`define LR_CONSTANT 0;
`define LR_ITER 1;
`define LR_DATA 2;
`define LR_HYBRID 3;
`define LR_DECAY LR_CONSTANT;
`define MAX_LEARNING_RATE 10;
`define BETA_LR 3;
`define RETRAIN 0;
`define VITIS_HLS_XILINX_PATH "C:/Xilinx/Vitis_HLS/2023.1/bin/vitis_hls.bat";
`define VIVADO_XILINX_PATH "C:/Xilinx/Vivado/2023.1/bin/vivado.bat";
`define VITIS_XILINX_PATH "C:/Xilinx/Vitis/2023.1/bin/vitis.bat";
