/**
 * @file level_hvec_gen_hdl.hpp
 * @brief This script generates HDL code for generating high-dimensional LEVEL vectors.
 * It is a novel method; for more information, please refer to our paper.
 *
 * @author Saeid Jamili and Marco Angioli
 * @note Author names are listed in alphabetical order.
 * @email <saeid.jamili@uniroma1.it>
 * @email <marco.angioli@uniroma1.it>
 *
 * @contributors
 *
 * @date Created: 24th July 2023
 * @date Last Updated: 23th August 2023
 *
 * @version 1.0.0
 *
 * @institute Sapienza University of Rome
 * @cite https://doi.org/10.xxxx/yyyyy
 *
 * @section DEPENDENCIES
 * - Dependency1: Description or version details.
 * - Dependency2: Description or version details.
 *
 * @section LICENSE
 * This file is part of the Aeneas HyperCompute Platform.
 *
 * Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 *
 * @section CHANGELOG
 * @version 1.0.0-dev - 23th August 2023
 * - Initial release
 *
 * @todo
 * - Complete level vector generator function
 * - Add training
 *
 * @see
 * -
 * -
 * -
 *
 */

module level_vec_gen (
    output reg [63:0] level_vec_out,
    input [2:0] frame_index,
    input [4:0] frame_id
);
    always @(*) begin
        // Update this function to match your requirements
        case (frame_index)
            0: begin
                case (frame_id)
                    0: level_vec_out = 64'b1010101110011010000001100011010101000001111011110100100001001001;
                    1: level_vec_out = 64'b1010101110111010000001100011010101000001111011110100100001001001;
                    2: level_vec_out = 64'b1010101110111010000001100111011101000001111011110100100001001001;
                    3: level_vec_out = 64'b1010101110111010000001100111011101000001111011110100100011001001;
                    4: level_vec_out = 64'b1010101110111010000001100111011101000001111011110100100011001001;
                    5: level_vec_out = 64'b1010101110111010000001100111011101000001111011110100100011001001;
                    6: level_vec_out = 64'b1010101110111010000001100111011101000001111011110100110011001001;
                    7: level_vec_out = 64'b1010101110111010000001100111011101000001111011110100110011001001;
                    8: level_vec_out = 64'b1010101110111010100001101111011101000001111011110101110011001001;
                    9: level_vec_out = 64'b1010101110111010100001101111011101000001111011110101110011001001;
                    10: level_vec_out = 64'b1110101110111010100001101111011101000001111011110101110011001001;
                    11: level_vec_out = 64'b1110101110111010100001101111011101001001111011110101110011001001;
                    12: level_vec_out = 64'b1110101110111010100001101111011101001011111011110101110011001001;
                    13: level_vec_out = 64'b1110101110111010100001101111011101001011111011110101110011001001;
                    14: level_vec_out = 64'b1110101110111010110001101111111101001011111011110101111011001001;
                    15: level_vec_out = 64'b1110101110111010110011101111111101001011111011110101111011001001;
                    16: level_vec_out = 64'b1110101110111010110011111111111101001011111011110101111011001001;
                    17: level_vec_out = 64'b1110101110111010110011111111111101001111111011110101111011001001;
                    18: level_vec_out = 64'b1111101110111010110011111111111101001111111011110101111011001001;
                    19: level_vec_out = 64'b1111101110111010110011111111111101001111111011110101111011101001;
                    20: level_vec_out = 64'b1111101110111110110011111111111101001111111011110101111011111001;
                    21: level_vec_out = 64'b1111101110111110110011111111111101001111111111110101111011111001;
                    22: level_vec_out = 64'b1111101110111110110011111111111101001111111111110101111011111001;
                    23: level_vec_out = 64'b1111101110111111110011111111111101001111111111110111111011111001;
                    24: level_vec_out = 64'b1111101110111111110011111111111101001111111111110111111011111001;
                    25: level_vec_out = 64'b1111101111111111110011111111111101001111111111110111111011111001;
                    26: level_vec_out = 64'b1111101111111111110011111111111101001111111111110111111011111001;
                    27: level_vec_out = 64'b1111101111111111111111111111111101101111111111110111111011111001;
                    28: level_vec_out = 64'b1111101111111111111111111111111101101111111111111111111011111101;
                    29: level_vec_out = 64'b1111101111111111111111111111111111101111111111111111111011111101;
                    30: level_vec_out = 64'b1111101111111111111111111111111111101111111111111111111011111101;
                    31: level_vec_out = 64'b1111101111111111111111111111111111111111111111111111111011111111;
                endcase
            end
            1: begin
                case (frame_id)
                    0: level_vec_out = 64'b0101000101111001100010111000001111001010001110010010111001001110;
                    1: level_vec_out = 64'b0101000101111001100010111000001111001010011110010010111001001110;
                    2: level_vec_out = 64'b0101000101111001100010111000001111001010011110010010111001001110;
                    3: level_vec_out = 64'b0101000101111001100010111010001111001010011111010010111001001110;
                    4: level_vec_out = 64'b0101000101111001100010111010001111001010011111010010111001001110;
                    5: level_vec_out = 64'b0101100101111001110010111010001111001010011111010010111001001110;
                    6: level_vec_out = 64'b0101100101111001110010111010001111001010011111110010111001001110;
                    7: level_vec_out = 64'b0101100101111001110010111010001111001010011111110010111001101111;
                    8: level_vec_out = 64'b0101100101111001110010111010001111001010011111110010111001101111;
                    9: level_vec_out = 64'b0101100101111001110110111010001111101010011111110010111001111111;
                    10: level_vec_out = 64'b0101100101111001110110111010001111101010011111110010111001111111;
                    11: level_vec_out = 64'b0101100101111001110110111010001111101010011111110010111001111111;
                    12: level_vec_out = 64'b0111100101111001110110111010001111101010011111110110111001111111;
                    13: level_vec_out = 64'b0111100101111001110110111010001111101011011111110110111101111111;
                    14: level_vec_out = 64'b0111100101111001110110111010001111101011011111110110111101111111;
                    15: level_vec_out = 64'b0111100101111001110110111010001111101011011111110110111101111111;
                    16: level_vec_out = 64'b0111110101111001110110111010011111101011011111110110111101111111;
                    17: level_vec_out = 64'b0111110101111001110110111010111111101011011111110110111101111111;
                    18: level_vec_out = 64'b0111110101111001110111111010111111101011011111110110111101111111;
                    19: level_vec_out = 64'b0111110101111001110111111010111111101011011111110110111101111111;
                    20: level_vec_out = 64'b0111110101111001110111111010111111101011011111110110111101111111;
                    21: level_vec_out = 64'b0111110101111011110111111010111111101011011111110110111101111111;
                    22: level_vec_out = 64'b0111111101111011111111111010111111101011011111110110111101111111;
                    23: level_vec_out = 64'b0111111101111111111111111010111111101011011111110110111111111111;
                    24: level_vec_out = 64'b1111111101111111111111111010111111101011011111110110111111111111;
                    25: level_vec_out = 64'b1111111101111111111111111010111111101011011111110110111111111111;
                    26: level_vec_out = 64'b1111111101111111111111111010111111111011011111110111111111111111;
                    27: level_vec_out = 64'b1111111111111111111111111010111111111111011111110111111111111111;
                    28: level_vec_out = 64'b1111111111111111111111111110111111111111011111110111111111111111;
                    29: level_vec_out = 64'b1111111111111111111111111110111111111111111111110111111111111111;
                    30: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    31: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                endcase
            end
            2: begin
                case (frame_id)
                    0: level_vec_out = 64'b1100110010010110001110110001110111010100111110101000100100010001;
                    1: level_vec_out = 64'b1100110010010110001110110001110111010100111110101000100100010001;
                    2: level_vec_out = 64'b1100110110010110001110110001110111010100111110101000100100010001;
                    3: level_vec_out = 64'b1100110110010110001110110001110111010100111110111010100100010001;
                    4: level_vec_out = 64'b1100110110010110001110110001110111010100111110111010100100010001;
                    5: level_vec_out = 64'b1100110110010110001110110011110111010110111110111010100100010001;
                    6: level_vec_out = 64'b1100110110010110001110110011110111110110111110111010101100010001;
                    7: level_vec_out = 64'b1101110110010110001110111011110111110110111110111010101100010001;
                    8: level_vec_out = 64'b1101110110010110001110111011110111110110111110111010101100010001;
                    9: level_vec_out = 64'b1101110110010110001110111011110111110110111110111010101100010001;
                    10: level_vec_out = 64'b1101110110010110001110111111110111110110111110111010101101010011;
                    11: level_vec_out = 64'b1111110110010110101110111111110111110110111110111110101101010011;
                    12: level_vec_out = 64'b1111110110010110101110111111110111110110111110111110101101010011;
                    13: level_vec_out = 64'b1111110110011110101110111111110111110110111110111110101101010011;
                    14: level_vec_out = 64'b1111110110011110101110111111110111110110111110111111101101110011;
                    15: level_vec_out = 64'b1111110110011110101110111111110111110110111110111111101101110011;
                    16: level_vec_out = 64'b1111110110011110101110111111110111110110111110111111101101110011;
                    17: level_vec_out = 64'b1111110110111110101110111111110111110110111110111111101101110011;
                    18: level_vec_out = 64'b1111110110111110101110111111110111110110111110111111101101111011;
                    19: level_vec_out = 64'b1111110110111110101110111111111111110111111110111111101111111011;
                    20: level_vec_out = 64'b1111110110111111111110111111111111110111111110111111101111111011;
                    21: level_vec_out = 64'b1111110110111111111110111111111111110111111110111111101111111011;
                    22: level_vec_out = 64'b1111110110111111111110111111111111110111111111111111111111111011;
                    23: level_vec_out = 64'b1111111110111111111111111111111111111111111111111111111111111011;
                    24: level_vec_out = 64'b1111111110111111111111111111111111111111111111111111111111111011;
                    25: level_vec_out = 64'b1111111110111111111111111111111111111111111111111111111111111011;
                    26: level_vec_out = 64'b1111111110111111111111111111111111111111111111111111111111111011;
                    27: level_vec_out = 64'b1111111110111111111111111111111111111111111111111111111111111011;
                    28: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111011;
                    29: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111011;
                    30: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111011;
                    31: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111011;
                endcase
            end
            3: begin
                case (frame_id)
                    0: level_vec_out = 64'b1101010011000100101111110011110110101101001001010001010010001100;
                    1: level_vec_out = 64'b1101010011000100101111110011110110101101101001010001010010001100;
                    2: level_vec_out = 64'b1101010011000100101111111011110110101101101001010001010010001100;
                    3: level_vec_out = 64'b1101010011000100101111111011110110101101101001010001010010001100;
                    4: level_vec_out = 64'b1101010011000100101111111011110110101101101001010001010010001101;
                    5: level_vec_out = 64'b1111010011000100101111111011110110101101101001010001010010001101;
                    6: level_vec_out = 64'b1111010011000100101111111011110110101101101001010001010010001101;
                    7: level_vec_out = 64'b1111010011010100101111111011110110101101101001010001010010001101;
                    8: level_vec_out = 64'b1111010011010100101111111011110110111101101001010001010010001101;
                    9: level_vec_out = 64'b1111010111010100101111111011110110111101101011010001010010001101;
                    10: level_vec_out = 64'b1111010111010100101111111011111110111101101011010001010010011101;
                    11: level_vec_out = 64'b1111010111010100101111111011111111111101101011010001010010011101;
                    12: level_vec_out = 64'b1111010111010100101111111011111111111101101011010001010110011101;
                    13: level_vec_out = 64'b1111010111010100101111111011111111111101101011010001010110011101;
                    14: level_vec_out = 64'b1111010111110110101111111011111111111101101011010001010110011101;
                    15: level_vec_out = 64'b1111010111110110101111111011111111111101101011010001010110011101;
                    16: level_vec_out = 64'b1111010111110110101111111011111111111101101011110001010110011101;
                    17: level_vec_out = 64'b1111010111110110101111111011111111111101101011110001010110011101;
                    18: level_vec_out = 64'b1111010111110110101111111011111111111111101011110001010110011101;
                    19: level_vec_out = 64'b1111010111110110101111111111111111111111101011110001010110011101;
                    20: level_vec_out = 64'b1111010111110110101111111111111111111111101011110001010110011101;
                    21: level_vec_out = 64'b1111010111110110111111111111111111111111101011110001010110011101;
                    22: level_vec_out = 64'b1111010111110111111111111111111111111111101011110101010110011101;
                    23: level_vec_out = 64'b1111010111110111111111111111111111111111101011110101010110011101;
                    24: level_vec_out = 64'b1111110111110111111111111111111111111111101011110111110110011101;
                    25: level_vec_out = 64'b1111110111110111111111111111111111111111101011110111111110011101;
                    26: level_vec_out = 64'b1111110111110111111111111111111111111111101111110111111110011101;
                    27: level_vec_out = 64'b1111110111110111111111111111111111111111101111110111111110011101;
                    28: level_vec_out = 64'b1111110111110111111111111111111111111111111111110111111110111101;
                    29: level_vec_out = 64'b1111111111110111111111111111111111111111111111110111111110111101;
                    30: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111110111101;
                    31: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111101;
                endcase
            end
            4: begin
                case (frame_id)
                    0: level_vec_out = 64'b1011100111100001100100010001101110110100000110111010000111111111;
                    1: level_vec_out = 64'b1011100111100001100100010001101110110100011110111010000111111111;
                    2: level_vec_out = 64'b1011100111110001100100010001101110111100011111111010000111111111;
                    3: level_vec_out = 64'b1011100111110001100100010001101110111100011111111010100111111111;
                    4: level_vec_out = 64'b1011100111110001100100010001101110111100011111111010100111111111;
                    5: level_vec_out = 64'b1011100111110001100100010001101110111100011111111010100111111111;
                    6: level_vec_out = 64'b1011100111110001100100010001101110111100011111111010100111111111;
                    7: level_vec_out = 64'b1011110111110001100100010001101110111100011111111010100111111111;
                    8: level_vec_out = 64'b1011110111110001100100010001101110111100111111111010100111111111;
                    9: level_vec_out = 64'b1011110111110001100100110001101110111101111111111010100111111111;
                    10: level_vec_out = 64'b1011110111110001100100110011101110111101111111111010100111111111;
                    11: level_vec_out = 64'b1011110111110001100100110011111110111101111111111010100111111111;
                    12: level_vec_out = 64'b1011110111110101100101110011111110111101111111111010100111111111;
                    13: level_vec_out = 64'b1011110111110101100101110011111110111101111111111010100111111111;
                    14: level_vec_out = 64'b1011110111110101100101110011111110111101111111111010100111111111;
                    15: level_vec_out = 64'b1011110111110101100101110011111110111101111111111010100111111111;
                    16: level_vec_out = 64'b1111110111110111100101110011111110111101111111111010100111111111;
                    17: level_vec_out = 64'b1111110111110111100101110011111110111101111111111010100111111111;
                    18: level_vec_out = 64'b1111110111110111100101110011111111111111111111111010100111111111;
                    19: level_vec_out = 64'b1111110111110111100101110011111111111111111111111010100111111111;
                    20: level_vec_out = 64'b1111110111110111100101110011111111111111111111111010100111111111;
                    21: level_vec_out = 64'b1111110111110111100101110011111111111111111111111110100111111111;
                    22: level_vec_out = 64'b1111110111110111100101110011111111111111111111111110101111111111;
                    23: level_vec_out = 64'b1111110111110111100101110011111111111111111111111110101111111111;
                    24: level_vec_out = 64'b1111110111110111101101110011111111111111111111111110101111111111;
                    25: level_vec_out = 64'b1111110111110111101101110011111111111111111111111110111111111111;
                    26: level_vec_out = 64'b1111111111111111111101110011111111111111111111111110111111111111;
                    27: level_vec_out = 64'b1111111111111111111101110011111111111111111111111110111111111111;
                    28: level_vec_out = 64'b1111111111111111111101111011111111111111111111111110111111111111;
                    29: level_vec_out = 64'b1111111111111111111111111011111111111111111111111110111111111111;
                    30: level_vec_out = 64'b1111111111111111111111111011111111111111111111111111111111111111;
                    31: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                endcase
            end
            5: begin
                case (frame_id)
                    0: level_vec_out = 64'b0000101001111100010010101011101110011001111100100101001100010110;
                    1: level_vec_out = 64'b0000101001111100010010101011101110011001111100100101011100010110;
                    2: level_vec_out = 64'b0000101001111100010010101011101110011001111100100101011100010110;
                    3: level_vec_out = 64'b0000101001111100010010101011101110011001111100100101011100010110;
                    4: level_vec_out = 64'b0000101001111100010011101011101110011001111101100101011100010110;
                    5: level_vec_out = 64'b0000101001111100010011101111101110011001111111100101011100010110;
                    6: level_vec_out = 64'b0000101001111100010011101111101110011001111111100101011100010110;
                    7: level_vec_out = 64'b0000101001111100010011101111101110011001111111100101011100010110;
                    8: level_vec_out = 64'b0000101001111100010111101111101110011001111111100101011100010110;
                    9: level_vec_out = 64'b0000101001111100010111101111101110011001111111100101011100010110;
                    10: level_vec_out = 64'b0000101001111100010111101111101110011001111111100101011100010110;
                    11: level_vec_out = 64'b0000101001111100010111101111101110011001111111100101011100010110;
                    12: level_vec_out = 64'b0000101001111100010111101111101110011001111111100101011100010110;
                    13: level_vec_out = 64'b0001101001111100010111101111101110011001111111100101111100010110;
                    14: level_vec_out = 64'b0001101001111100010111101111101110011001111111100101111100010110;
                    15: level_vec_out = 64'b0101101001111100010111111111101110011001111111100101111100010110;
                    16: level_vec_out = 64'b0111101001111100010111111111101110011001111111100101111100010110;
                    17: level_vec_out = 64'b0111111001111100010111111111101110011001111111100111111100010110;
                    18: level_vec_out = 64'b0111111001111100011111111111101110111001111111100111111100010110;
                    19: level_vec_out = 64'b0111111001111100011111111111101111111001111111100111111100010110;
                    20: level_vec_out = 64'b0111111001111110011111111111111111111001111111100111111100010110;
                    21: level_vec_out = 64'b0111111011111110011111111111111111111001111111100111111100010110;
                    22: level_vec_out = 64'b0111111011111110011111111111111111111001111111100111111100010110;
                    23: level_vec_out = 64'b0111111011111110011111111111111111111001111111110111111100010110;
                    24: level_vec_out = 64'b0111111011111110011111111111111111111001111111110111111100011111;
                    25: level_vec_out = 64'b1111111111111110011111111111111111111101111111110111111100011111;
                    26: level_vec_out = 64'b1111111111111110011111111111111111111101111111110111111110011111;
                    27: level_vec_out = 64'b1111111111111110011111111111111111111101111111110111111110111111;
                    28: level_vec_out = 64'b1111111111111110011111111111111111111101111111110111111110111111;
                    29: level_vec_out = 64'b1111111111111110011111111111111111111101111111111111111110111111;
                    30: level_vec_out = 64'b1111111111111111011111111111111111111101111111111111111110111111;
                    31: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111110111111;
                endcase
            end
            6: begin
                case (frame_id)
                    0: level_vec_out = 64'b0011000110001011001010010111100001011011110010111110000001011010;
                    1: level_vec_out = 64'b0111000110001011001010011111100001011011110010111110000001011010;
                    2: level_vec_out = 64'b0111000110001011001010011111100001011011110010111110000001011010;
                    3: level_vec_out = 64'b0111000110001011001010011111100001011011110010111110000001011010;
                    4: level_vec_out = 64'b0111000110001011001010011111100001011011110010111110000001011011;
                    5: level_vec_out = 64'b0111001110001011001010011111100001011011110010111110000001011011;
                    6: level_vec_out = 64'b0111101110001011001010111111100001011011110011111110000001011011;
                    7: level_vec_out = 64'b0111101110001011001010111111100001011011110011111110000001011111;
                    8: level_vec_out = 64'b0111101110001011001010111111100001011011110011111111000001011111;
                    9: level_vec_out = 64'b0111101110001011001010111111100001011011110011111111000001011111;
                    10: level_vec_out = 64'b0111101110101011001010111111100001011011110011111111000001011111;
                    11: level_vec_out = 64'b0111101110101011001010111111100011011111110011111111000001011111;
                    12: level_vec_out = 64'b0111101110101011001010111111100011011111110011111111000111011111;
                    13: level_vec_out = 64'b0111101110101011001010111111100011011111110011111111100111011111;
                    14: level_vec_out = 64'b0111101110101011001010111111100011011111110011111111100111011111;
                    15: level_vec_out = 64'b0111101110111011001010111111100011011111111011111111100111011111;
                    16: level_vec_out = 64'b0111101110111011001010111111100011011111111111111111100111011111;
                    17: level_vec_out = 64'b0111101110111011001010111111100111011111111111111111100111011111;
                    18: level_vec_out = 64'b0111101110111011001010111111100111011111111111111111100111011111;
                    19: level_vec_out = 64'b0111101110111011001010111111100111111111111111111111100111011111;
                    20: level_vec_out = 64'b0111101110111011001010111111100111111111111111111111100111011111;
                    21: level_vec_out = 64'b0111101110111011001010111111111111111111111111111111100111011111;
                    22: level_vec_out = 64'b0111101110111011001010111111111111111111111111111111100111011111;
                    23: level_vec_out = 64'b0111101110111011001010111111111111111111111111111111100111011111;
                    24: level_vec_out = 64'b0111101110111011011010111111111111111111111111111111100111011111;
                    25: level_vec_out = 64'b0111101110111011011011111111111111111111111111111111100111111111;
                    26: level_vec_out = 64'b0111101110111011011011111111111111111111111111111111100111111111;
                    27: level_vec_out = 64'b0111101111111011011011111111111111111111111111111111110111111111;
                    28: level_vec_out = 64'b0111101111111011011111111111111111111111111111111111110111111111;
                    29: level_vec_out = 64'b1111101111111011011111111111111111111111111111111111110111111111;
                    30: level_vec_out = 64'b1111101111111111011111111111111111111111111111111111111111111111;
                    31: level_vec_out = 64'b1111101111111111011111111111111111111111111111111111111111111111;
                endcase
            end
            7: begin
                case (frame_id)
                    0: level_vec_out = 64'b0000111011010011101110100100010011100001101100111101111101000110;
                    1: level_vec_out = 64'b0000111011010011101110100100010011100001101100111101111101000110;
                    2: level_vec_out = 64'b0000111011011011101110100100010011100001101100111101111101000110;
                    3: level_vec_out = 64'b0000111011011011101110110100011011100001101100111101111101000110;
                    4: level_vec_out = 64'b0001111011011011101110110110011011100001101100111101111111001110;
                    5: level_vec_out = 64'b0001111011011011101110110110011011100001101100111101111111001110;
                    6: level_vec_out = 64'b0001111011011011101110110110011011100001101100111101111111011110;
                    7: level_vec_out = 64'b0001111011011011101110110110011011100001101101111101111111011110;
                    8: level_vec_out = 64'b0011111011011011101110110110011011100001101101111101111111011110;
                    9: level_vec_out = 64'b0111111011011011101110110110011011100001101101111101111111011110;
                    10: level_vec_out = 64'b0111111011011011101110110110011011100001101101111101111111011110;
                    11: level_vec_out = 64'b0111111011011011101110110110011011100001101101111101111111011110;
                    12: level_vec_out = 64'b0111111011011011101110110110011011100001101101111101111111011110;
                    13: level_vec_out = 64'b0111111011011011101110110110011011110001101101111101111111111110;
                    14: level_vec_out = 64'b0111111011011011101110110110011011110001111101111101111111111110;
                    15: level_vec_out = 64'b1111111011011011101111110111011011110001111101111101111111111110;
                    16: level_vec_out = 64'b1111111011011011101111110111011011110001111101111101111111111110;
                    17: level_vec_out = 64'b1111111011011011101111110111011011110011111101111101111111111111;
                    18: level_vec_out = 64'b1111111011011011101111110111011011110011111101111101111111111111;
                    19: level_vec_out = 64'b1111111011011011101111110111111011110011111101111101111111111111;
                    20: level_vec_out = 64'b1111111011011011101111110111111011111011111111111101111111111111;
                    21: level_vec_out = 64'b1111111011111011101111110111111011111011111111111101111111111111;
                    22: level_vec_out = 64'b1111111011111011101111110111111111111011111111111101111111111111;
                    23: level_vec_out = 64'b1111111011111011101111110111111111111011111111111101111111111111;
                    24: level_vec_out = 64'b1111111011111011101111110111111111111011111111111101111111111111;
                    25: level_vec_out = 64'b1111111011111011101111110111111111111011111111111101111111111111;
                    26: level_vec_out = 64'b1111111011111111101111110111111111111011111111111101111111111111;
                    27: level_vec_out = 64'b1111111011111111101111110111111111111011111111111101111111111111;
                    28: level_vec_out = 64'b1111111011111111101111110111111111111011111111111101111111111111;
                    29: level_vec_out = 64'b1111111011111111111111110111111111111011111111111111111111111111;
                    30: level_vec_out = 64'b1111111011111111111111110111111111111011111111111111111111111111;
                    31: level_vec_out = 64'b1111111111111111111111110111111111111111111111111111111111111111;
                endcase
            end
        endcase
    end
endmodule