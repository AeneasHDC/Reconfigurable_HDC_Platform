----
 -- @file level_hvec_gen_hdl.hpp
 -- @brief This script generates HDL code for generating high-dimensional LEVEL vectors.
 -- It is a novel method; for more information, please refer to our paper.
 --
 -- @author Saeid Jamili and Marco Angioli
 -- @note Author names are listed in alphabetical order.
 -- @email <saeid.jamili@uniroma1.it>
 -- @email <marco.angioli@uniroma1.it>
 --
 -- @contributors
 --
 -- @date Created: 24th July 2023
 -- @date Last Updated: 23th August 2023
 --
 -- @version 1.0.0
 --
 -- @institute Sapienza University of Rome
 -- @cite https://doi.org/10.xxxx/yyyyy
 --
 -- @section DEPENDENCIES
 -- - Dependency1: Description or version details.
 -- - Dependency2: Description or version details.
 --
 -- @section LICENSE
 -- This file is part of the Aeneas HyperCompute Platform.
 --
 -- Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 --
 -- @section CHANGELOG
 -- @version 1.0.0-dev - 23th August 2023
 -- - Initial release
 --
 -- @todo
 -- - Complete level vector generator function
 -- - Add training
 --
 -- @see
 -- -
 -- -
 -- -
 --
 --

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity level_vec_gen is
    Port ( level_vec_out : out  STD_LOGIC_VECTOR (63 downto 0);
           frame_index : in  STD_LOGIC_VECTOR (2 downto 0);
           frame_id : in  STD_LOGIC_VECTOR (4 downto 0));
end level_vec_gen;

architecture Behavioral of level_vec_gen is
begin
    process (frame_index, frame_id)
    begin
        -- Update this function to match your requirements
        case frame_index is
            when "000" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0100110001000111011001110111101011000110100010010000100110100101";
                    when "00001" => level_vec_out <= "0100110001000111011001110111101011000110110010010000100110100101";
                    when "00010" => level_vec_out <= "0100110001000111011001111111101011000110110010010000100110100101";
                    when "00011" => level_vec_out <= "0100111001000111011011111111101011000110110010010000110110100101";
                    when "00100" => level_vec_out <= "0100111001000111011011111111101011000110110010110000110110100101";
                    when "00101" => level_vec_out <= "0100111001100111011011111111101011000110110010110100110110100101";
                    when "00110" => level_vec_out <= "0100111001100111011011111111101011000110110011110110110110100101";
                    when "00111" => level_vec_out <= "0100111001100111011011111111101011000110110011110110110110100101";
                    when "01000" => level_vec_out <= "0101111001100111011011111111101011000110110011110110110110100101";
                    when "01001" => level_vec_out <= "0101111001100111011011111111101011000110110011110110110110100101";
                    when "01010" => level_vec_out <= "1101111011100111011011111111101011000110110011110110110110100101";
                    when "01011" => level_vec_out <= "1101111011101111011111111111101011000110110011110110110110101101";
                    when "01100" => level_vec_out <= "1101111011101111011111111111101011000110110011110110110110101101";
                    when "01101" => level_vec_out <= "1101111011111111011111111111101011000110110011110110111110101101";
                    when "01110" => level_vec_out <= "1101111011111111011111111111101111000110110011110110111110101101";
                    when "01111" => level_vec_out <= "1101111011111111011111111111101111000110111011110110111110101101";
                    when "10000" => level_vec_out <= "1101111011111111011111111111101111000110111011110110111110101101";
                    when "10001" => level_vec_out <= "1101111011111111011111111111101111000110111011110110111110101101";
                    when "10010" => level_vec_out <= "1101111011111111011111111111101111000110111011110111111110101101";
                    when "10011" => level_vec_out <= "1101111011111111011111111111101111000110111011110111111110101101";
                    when "10100" => level_vec_out <= "1101111011111111011111111111101111000111111011110111111110101101";
                    when "10101" => level_vec_out <= "1101111011111111011111111111111111000111111011110111111110101101";
                    when "10110" => level_vec_out <= "1101111011111111011111111111111111000111111011110111111110101101";
                    when "10111" => level_vec_out <= "1101111011111111011111111111111111000111111011110111111110101101";
                    when "11000" => level_vec_out <= "1101111011111111011111111111111111110111111011110111111110111101";
                    when "11001" => level_vec_out <= "1101111011111111011111111111111111110111111011110111111110111101";
                    when "11010" => level_vec_out <= "1111111011111111111111111111111111110111111011110111111111111101";
                    when "11011" => level_vec_out <= "1111111011111111111111111111111111110111111111110111111111111111";
                    when "11100" => level_vec_out <= "1111111011111111111111111111111111110111111111110111111111111111";
                    when "11101" => level_vec_out <= "1111111011111111111111111111111111110111111111110111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111110111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111110111111111111111111111111111";
                when others => null;
                end case;
            when "001" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1101000100101100101000010011100100100101101000111010100101001000";
                    when "00001" => level_vec_out <= "1101000100101100101000010011100100100101101000111010100101001000";
                    when "00010" => level_vec_out <= "1111000100101100101000010011100100100101101000111010100101001000";
                    when "00011" => level_vec_out <= "1111000100101100101000010011100100100101101000111010100101001000";
                    when "00100" => level_vec_out <= "1111000100101100101000010011100100100101101000111010100101001000";
                    when "00101" => level_vec_out <= "1111000110101100101000011011100100100101101000111010100101001000";
                    when "00110" => level_vec_out <= "1111100110101100101000011011100100100101101001111010100101001000";
                    when "00111" => level_vec_out <= "1111100110101100101000011011100100100101101011111010100101001000";
                    when "01000" => level_vec_out <= "1111100110101100101000011011100100100101101011111010100101001000";
                    when "01001" => level_vec_out <= "1111100110101100101000011011100100100101101111111010100101001000";
                    when "01010" => level_vec_out <= "1111100110101100101100011011100100100101101111111010100101001000";
                    when "01011" => level_vec_out <= "1111100110101100101100011011100100100101101111111010100101001000";
                    when "01100" => level_vec_out <= "1111100110101110101100011011100100100101111111111010100101001000";
                    when "01101" => level_vec_out <= "1111100110101110101100011011100100100101111111111010100101001000";
                    when "01110" => level_vec_out <= "1111100111101110101100111011100100100101111111111010100101001000";
                    when "01111" => level_vec_out <= "1111100111101110101101111011110100100101111111111010100101001000";
                    when "10000" => level_vec_out <= "1111100111101110101101111011110100100101111111111010100101001000";
                    when "10001" => level_vec_out <= "1111100111101110101101111011110100100101111111111010100101001000";
                    when "10010" => level_vec_out <= "1111100111101111101101111011110100100111111111111110100111001000";
                    when "10011" => level_vec_out <= "1111100111101111101101111011110100100111111111111110101111001000";
                    when "10100" => level_vec_out <= "1111100111101111101101111011110100100111111111111110101111001100";
                    when "10101" => level_vec_out <= "1111100111101111101101111011110110100111111111111110101111001100";
                    when "10110" => level_vec_out <= "1111110111101111101101111011111110100111111111111110101111001100";
                    when "10111" => level_vec_out <= "1111110111101111101101111011111111100111111111111110101111001100";
                    when "11000" => level_vec_out <= "1111110111101111101101111011111111100111111111111110101111001100";
                    when "11001" => level_vec_out <= "1111111111101111101101111011111111110111111111111110101111011100";
                    when "11010" => level_vec_out <= "1111111111101111101101111011111111110111111111111110101111011100";
                    when "11011" => level_vec_out <= "1111111111101111101101111011111111110111111111111111101111011100";
                    when "11100" => level_vec_out <= "1111111111111111101101111011111111110111111111111111101111111110";
                    when "11101" => level_vec_out <= "1111111111111111101111111011111111111111111111111111101111111110";
                    when "11110" => level_vec_out <= "1111111111111111101111111111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111101111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "010" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1001011000101111001100110111010000001101010000000001000110001101";
                    when "00001" => level_vec_out <= "1001011000101111001100110111010000001101010100000001000110001101";
                    when "00010" => level_vec_out <= "1001011000101111001110110111011000001101010100000001000110001101";
                    when "00011" => level_vec_out <= "1001011000101111001110110111011000001101010100000001000110001111";
                    when "00100" => level_vec_out <= "1001011000101111001110110111011000001101010100000001000110001111";
                    when "00101" => level_vec_out <= "1001011100101111001110110111011001001101010100000001000110001111";
                    when "00110" => level_vec_out <= "1001011100101111001110110111011001001101010100000001000110001111";
                    when "00111" => level_vec_out <= "1001011100101111001110111111011001001101010100000001000110001111";
                    when "01000" => level_vec_out <= "1001011100101111101110111111011011001101010100000001000110001111";
                    when "01001" => level_vec_out <= "1001011100101111101110111111011011001101010100000001000110001111";
                    when "01010" => level_vec_out <= "1001011100111111101110111111011011001101010100000001000110001111";
                    when "01011" => level_vec_out <= "1001011110111111101110111111011111001101010100000001000110001111";
                    when "01100" => level_vec_out <= "1001011110111111111110111111011111001101010100000001000111001111";
                    when "01101" => level_vec_out <= "1001011110111111111111111111011111001101010100000011000111001111";
                    when "01110" => level_vec_out <= "1001111110111111111111111111011111001111010100000011010111001111";
                    when "01111" => level_vec_out <= "1001111110111111111111111111011111001111010100000011010111001111";
                    when "10000" => level_vec_out <= "1001111110111111111111111111011111001111010110000011010111001111";
                    when "10001" => level_vec_out <= "1001111110111111111111111111011111001111010110000011010111101111";
                    when "10010" => level_vec_out <= "1001111110111111111111111111011111001111010111000011010111101111";
                    when "10011" => level_vec_out <= "1001111110111111111111111111011111001111010111000011010111101111";
                    when "10100" => level_vec_out <= "1001111110111111111111111111011111101111010111001011010111111111";
                    when "10101" => level_vec_out <= "1001111110111111111111111111011111101111010111001011010111111111";
                    when "10110" => level_vec_out <= "1011111110111111111111111111011111101111110111001011010111111111";
                    when "10111" => level_vec_out <= "1011111110111111111111111111011111101111110111001011011111111111";
                    when "11000" => level_vec_out <= "1011111110111111111111111111011111101111111111001011011111111111";
                    when "11001" => level_vec_out <= "1011111110111111111111111111011111111111111111001111011111111111";
                    when "11010" => level_vec_out <= "1011111110111111111111111111011111111111111111001111011111111111";
                    when "11011" => level_vec_out <= "1011111110111111111111111111011111111111111111001111011111111111";
                    when "11100" => level_vec_out <= "1111111110111111111111111111011111111111111111001111011111111111";
                    when "11101" => level_vec_out <= "1111111110111111111111111111011111111111111111111111011111111111";
                    when "11110" => level_vec_out <= "1111111110111111111111111111011111111111111111111111011111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111011111111111111111111111011111111111";
                when others => null;
                end case;
            when "011" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0100110001001010000000000101100111011010010011000110010100001111";
                    when "00001" => level_vec_out <= "0100110001001010000000000101100111011010010111000110010100001111";
                    when "00010" => level_vec_out <= "0100110001011010000000000101100111011010010111000110010100001111";
                    when "00011" => level_vec_out <= "0100110001011010000000000101100111011010010111000110010110001111";
                    when "00100" => level_vec_out <= "0100110001011010000000000101100111011010010111000110010110001111";
                    when "00101" => level_vec_out <= "0100110001011010000000000101100111011010010111010110010110001111";
                    when "00110" => level_vec_out <= "0100110101011010000000000101100111011010010111010110010110001111";
                    when "00111" => level_vec_out <= "0100110101011110000000000101100111011010011111010110010110001111";
                    when "01000" => level_vec_out <= "0100110101011110000100000101100111011011011111010110010110001111";
                    when "01001" => level_vec_out <= "0100110101011110000101000101100111011011011111010110010110011111";
                    when "01010" => level_vec_out <= "0100110101011110000101000101100111011011011111010110110110011111";
                    when "01011" => level_vec_out <= "0100110111011110000101000101100111011011011111010110110110011111";
                    when "01100" => level_vec_out <= "0100110111111110000101000101100111011011011111010110110110011111";
                    when "01101" => level_vec_out <= "0100110111111110000101000101100111011011011111011110110110011111";
                    when "01110" => level_vec_out <= "0100110111111110000101000101100111011011011111011110110110011111";
                    when "01111" => level_vec_out <= "0100110111111110010101000101100111111011011111011110110110011111";
                    when "10000" => level_vec_out <= "0100110111111110010101000101100111111011011111111110110110011111";
                    when "10001" => level_vec_out <= "1100110111111110010101100101100111111011011111111110110111011111";
                    when "10010" => level_vec_out <= "1100110111111110010101110101100111111011011111111110110111011111";
                    when "10011" => level_vec_out <= "1100110111111110010111110101100111111011111111111111110111011111";
                    when "10100" => level_vec_out <= "1100111111111110010111110101100111111011111111111111110111011111";
                    when "10101" => level_vec_out <= "1110111111111110010111110101100111111011111111111111110111011111";
                    when "10110" => level_vec_out <= "1110111111111110010111110101110111111011111111111111110111011111";
                    when "10111" => level_vec_out <= "1110111111111110010111110101110111111011111111111111110111111111";
                    when "11000" => level_vec_out <= "1110111111111111010111110101110111111011111111111111110111111111";
                    when "11001" => level_vec_out <= "1110111111111111110111110101110111111011111111111111110111111111";
                    when "11010" => level_vec_out <= "1110111111111111110111110111110111111111111111111111110111111111";
                    when "11011" => level_vec_out <= "1111111111111111110111111111110111111111111111111111111111111111";
                    when "11100" => level_vec_out <= "1111111111111111110111111111110111111111111111111111111111111111";
                    when "11101" => level_vec_out <= "1111111111111111111111111111110111111111111111111111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111110111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "100" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1110011000111001011110111000000011110001110101000101010011010101";
                    when "00001" => level_vec_out <= "1110011000111001011110111000000011110001110101000101010111010101";
                    when "00010" => level_vec_out <= "1110011000111001011110111000000011110001110101000101010111010101";
                    when "00011" => level_vec_out <= "1110011010111001011110111000000011110001110101000101010111010101";
                    when "00100" => level_vec_out <= "1110011010111101011110111000000011110001110101000101010111011101";
                    when "00101" => level_vec_out <= "1110011010111101011110111000000011110001110101000101010111011101";
                    when "00110" => level_vec_out <= "1110011010111101011110111000000011110001110101000101010111011101";
                    when "00111" => level_vec_out <= "1110011010111101011110111000000011110001110101000101010111011111";
                    when "01000" => level_vec_out <= "1111111010111101011110111010000011110001110101000101010111011111";
                    when "01001" => level_vec_out <= "1111111010111101111110111010000011110001110101000101010111111111";
                    when "01010" => level_vec_out <= "1111111010111101111110111010000011110001110101000101010111111111";
                    when "01011" => level_vec_out <= "1111111010111101111110111011000011110001110101000101010111111111";
                    when "01100" => level_vec_out <= "1111111010111111111110111011000011110001110101000101010111111111";
                    when "01101" => level_vec_out <= "1111111010111111111110111011000011110001110101010101010111111111";
                    when "01110" => level_vec_out <= "1111111011111111111110111011000011110001110101010101010111111111";
                    when "01111" => level_vec_out <= "1111111011111111111110111011000011111001110101010111010111111111";
                    when "10000" => level_vec_out <= "1111111011111111111110111011000011111001110101010111010111111111";
                    when "10001" => level_vec_out <= "1111111011111111111110111011001011111001110101010111010111111111";
                    when "10010" => level_vec_out <= "1111111011111111111111111011001011111001110101010111010111111111";
                    when "10011" => level_vec_out <= "1111111011111111111111111011001011111001110101010111010111111111";
                    when "10100" => level_vec_out <= "1111111111111111111111111011001011111001110101010111010111111111";
                    when "10101" => level_vec_out <= "1111111111111111111111111011011011111011110101010111010111111111";
                    when "10110" => level_vec_out <= "1111111111111111111111111011011011111011110111010111010111111111";
                    when "10111" => level_vec_out <= "1111111111111111111111111111011011111011110111010111111111111111";
                    when "11000" => level_vec_out <= "1111111111111111111111111111011111111011110111010111111111111111";
                    when "11001" => level_vec_out <= "1111111111111111111111111111011111111011110111010111111111111111";
                    when "11010" => level_vec_out <= "1111111111111111111111111111011111111011110111010111111111111111";
                    when "11011" => level_vec_out <= "1111111111111111111111111111011111111011110111010111111111111111";
                    when "11100" => level_vec_out <= "1111111111111111111111111111011111111111110111011111111111111111";
                    when "11101" => level_vec_out <= "1111111111111111111111111111011111111111110111111111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111011111111111110111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111110111111111111111111111";
                when others => null;
                end case;
            when "101" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0101110101111000111011011101010011110110111001111101010111010000";
                    when "00001" => level_vec_out <= "0101110101111000111011011101010011110110111001111101010111010000";
                    when "00010" => level_vec_out <= "0101110101111000111011011101011011110110111001111101010111010000";
                    when "00011" => level_vec_out <= "0101110101111000111011011101011011110110111001111111110111010000";
                    when "00100" => level_vec_out <= "0101110111111000111011011101011011110110111001111111110111110000";
                    when "00101" => level_vec_out <= "0101110111111000111011011101011011110110111001111111110111110000";
                    when "00110" => level_vec_out <= "0101110111111000111011011101011011110110111001111111110111110010";
                    when "00111" => level_vec_out <= "0101110111111000111011011101011011110110111001111111111111110010";
                    when "01000" => level_vec_out <= "0101110111111000111011011101011011110110111001111111111111110010";
                    when "01001" => level_vec_out <= "0101110111111000111011011101011011110111111001111111111111110010";
                    when "01010" => level_vec_out <= "0101110111111000111011011101011011110111111001111111111111110010";
                    when "01011" => level_vec_out <= "0101110111111000111011011101011011110111111001111111111111110010";
                    when "01100" => level_vec_out <= "0101110111111000111011011101011011111111111001111111111111110010";
                    when "01101" => level_vec_out <= "0101110111111001111011011101011011111111111001111111111111111010";
                    when "01110" => level_vec_out <= "0101110111111001111011111101011011111111111001111111111111111010";
                    when "01111" => level_vec_out <= "0101110111111001111011111101011011111111111001111111111111111010";
                    when "10000" => level_vec_out <= "0101110111111101111011111101011011111111111001111111111111111011";
                    when "10001" => level_vec_out <= "0101110111111101111011111101011011111111111101111111111111111111";
                    when "10010" => level_vec_out <= "0101110111111101111011111101011011111111111101111111111111111111";
                    when "10011" => level_vec_out <= "0101110111111101111011111111011011111111111101111111111111111111";
                    when "10100" => level_vec_out <= "0101110111111101111011111111011011111111111111111111111111111111";
                    when "10101" => level_vec_out <= "0101110111111101111011111111011011111111111111111111111111111111";
                    when "10110" => level_vec_out <= "0101110111111101111011111111011011111111111111111111111111111111";
                    when "10111" => level_vec_out <= "0111110111111101111011111111011011111111111111111111111111111111";
                    when "11000" => level_vec_out <= "0111110111111101111111111111011011111111111111111111111111111111";
                    when "11001" => level_vec_out <= "0111110111111111111111111111011011111111111111111111111111111111";
                    when "11010" => level_vec_out <= "1111110111111111111111111111011011111111111111111111111111111111";
                    when "11011" => level_vec_out <= "1111110111111111111111111111011011111111111111111111111111111111";
                    when "11100" => level_vec_out <= "1111110111111111111111111111111011111111111111111111111111111111";
                    when "11101" => level_vec_out <= "1111110111111111111111111111111111111111111111111111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "110" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0111011001100000011011100111110010011100100110101101111000100001";
                    when "00001" => level_vec_out <= "0111011001100001011011100111110010111100101111101101111000100001";
                    when "00010" => level_vec_out <= "0111011001100001011011100111110010111100101111101111111000100001";
                    when "00011" => level_vec_out <= "0111011001100001011011100111110010111100101111101111111000100001";
                    when "00100" => level_vec_out <= "0111011001100001011011100111110010111100101111101111111001100001";
                    when "00101" => level_vec_out <= "0111011001100001011011100111110010111100101111101111111001110001";
                    when "00110" => level_vec_out <= "0111011001100001011011100111110010111100101111101111111001110101";
                    when "00111" => level_vec_out <= "0111011001100001011011100111110010111100101111101111111001110101";
                    when "01000" => level_vec_out <= "0111011001100001011011100111110010111100101111101111111001110101";
                    when "01001" => level_vec_out <= "0111011001100001011011100111110010111100101111101111111011110101";
                    when "01010" => level_vec_out <= "0111011001100001011111100111110011111101101111101111111011110101";
                    when "01011" => level_vec_out <= "0111011001100001111111100111110011111101101111101111111011110101";
                    when "01100" => level_vec_out <= "0111011001100001111111100111111011111101101111101111111011110101";
                    when "01101" => level_vec_out <= "0111011001100001111111100111111011111101101111101111111011110101";
                    when "01110" => level_vec_out <= "0111011001100001111111100111111011111101101111101111111011110101";
                    when "01111" => level_vec_out <= "0111011001100101111111100111111011111101101111101111111011110101";
                    when "10000" => level_vec_out <= "0111111011100101111111100111111011111101101111101111111111110101";
                    when "10001" => level_vec_out <= "0111111011100101111111101111111011111101101111101111111111110101";
                    when "10010" => level_vec_out <= "0111111011100101111111101111111011111101101111101111111111110101";
                    when "10011" => level_vec_out <= "0111111011100101111111101111111011111101101111101111111111110101";
                    when "10100" => level_vec_out <= "0111111011100101111111101111111011111101101111101111111111110101";
                    when "10101" => level_vec_out <= "0111111011100101111111101111111111111111101111101111111111110101";
                    when "10110" => level_vec_out <= "0111111011100101111111101111111111111111101111101111111111110101";
                    when "10111" => level_vec_out <= "0111111011100101111111101111111111111111111111101111111111110101";
                    when "11000" => level_vec_out <= "0111111011100101111111101111111111111111111111101111111111110101";
                    when "11001" => level_vec_out <= "0111111111100101111111101111111111111111111111101111111111110101";
                    when "11010" => level_vec_out <= "0111111111100101111111101111111111111111111111101111111111110101";
                    when "11011" => level_vec_out <= "0111111111110101111111101111111111111111111111101111111111110101";
                    when "11100" => level_vec_out <= "0111111111110101111111101111111111111111111111101111111111110101";
                    when "11101" => level_vec_out <= "0111111111110101111111101111111111111111111111101111111111110101";
                    when "11110" => level_vec_out <= "0111111111110101111111101111111111111111111111101111111111111101";
                    when "11111" => level_vec_out <= "1111111111111101111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "111" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0010011101110101111111111101101000111101011100101110010101011110";
                    when "00001" => level_vec_out <= "0010011101110101111111111101101000111101011100101110010101011110";
                    when "00010" => level_vec_out <= "0010011101111101111111111101101000111101011100101110010101011110";
                    when "00011" => level_vec_out <= "0010011101111101111111111101101000111101011100101110010101011110";
                    when "00100" => level_vec_out <= "0010011101111101111111111101101000111111011100101110110101011110";
                    when "00101" => level_vec_out <= "0010011101111101111111111101101000111111011100101110110101011110";
                    when "00110" => level_vec_out <= "0010011101111101111111111101101000111111111100101110110101011110";
                    when "00111" => level_vec_out <= "0010011101111101111111111101101010111111111100111110110101011110";
                    when "01000" => level_vec_out <= "0010011101111101111111111101101010111111111100111110110101011110";
                    when "01001" => level_vec_out <= "0010011101111101111111111101101010111111111100111110111101011110";
                    when "01010" => level_vec_out <= "0010011101111101111111111101101010111111111100111110111101011110";
                    when "01011" => level_vec_out <= "0010011101111101111111111101101010111111111100111110111101011110";
                    when "01100" => level_vec_out <= "0010011101111101111111111101101010111111111100111110111101011110";
                    when "01101" => level_vec_out <= "0010011101111101111111111101101010111111111100111110111101011110";
                    when "01110" => level_vec_out <= "0010011101111101111111111101101010111111111100111110111101011110";
                    when "01111" => level_vec_out <= "0010011101111101111111111101101010111111111100111110111101011110";
                    when "10000" => level_vec_out <= "0011011101111101111111111101101010111111111100111110111101011110";
                    when "10001" => level_vec_out <= "0011011101111101111111111101101010111111111100111110111101011110";
                    when "10010" => level_vec_out <= "0011011101111101111111111101101010111111111100111110111101011110";
                    when "10011" => level_vec_out <= "0011011101111101111111111111101011111111111100111111111101011110";
                    when "10100" => level_vec_out <= "0011011101111101111111111111101011111111111100111111111101011110";
                    when "10101" => level_vec_out <= "0011011101111111111111111111101011111111111100111111111101011110";
                    when "10110" => level_vec_out <= "0011111101111111111111111111101011111111111100111111111111011110";
                    when "10111" => level_vec_out <= "0011111101111111111111111111101011111111111100111111111111011110";
                    when "11000" => level_vec_out <= "0111111101111111111111111111101011111111111100111111111111011110";
                    when "11001" => level_vec_out <= "0111111101111111111111111111101011111111111100111111111111011110";
                    when "11010" => level_vec_out <= "0111111101111111111111111111111011111111111100111111111111011111";
                    when "11011" => level_vec_out <= "1111111101111111111111111111111011111111111100111111111111011111";
                    when "11100" => level_vec_out <= "1111111111111111111111111111111011111111111100111111111111011111";
                    when "11101" => level_vec_out <= "1111111111111111111111111111111011111111111100111111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111011111111111101111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111011111111111101111111111111111111";
                when others => null;
                end case;
            when others => null;
        end case;
    end process;
end Behavioral;