----
 -- @file level_hvec_gen_hdl.hpp
 -- @brief This script generates HDL code for generating high-dimensional LEVEL vectors.
 -- It is a novel method; for more information, please refer to our paper.
 --
 -- @author Saeid Jamili and Marco Angioli
 -- @note Author names are listed in alphabetical order.
 -- @email <saeid.jamili@uniroma1.it>
 -- @email <marco.angioli@uniroma1.it>
 --
 -- @contributors
 --
 -- @date Created: 24th July 2023
 -- @date Last Updated: 23th August 2023
 --
 -- @version 1.0.0
 --
 -- @institute Sapienza University of Rome
 -- @cite https://doi.org/10.xxxx/yyyyy
 --
 -- @section DEPENDENCIES
 -- - Dependency1: Description or version details.
 -- - Dependency2: Description or version details.
 --
 -- @section LICENSE
 -- This file is part of the Aeneas HyperCompute Platform.
 --
 -- Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 --
 -- @section CHANGELOG
 -- @version 1.0.0-dev - 23th August 2023
 -- - Initial release
 --
 -- @todo
 -- - Complete level vector generator function
 -- - Add training
 --
 -- @see
 -- -
 -- -
 -- -
 --
 --

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity level_vec_gen is
    Port ( level_vec_out : out  STD_LOGIC_VECTOR (63 downto 0);
           frame_index : in  STD_LOGIC_VECTOR (2 downto 0);
           frame_id : in  STD_LOGIC_VECTOR (4 downto 0));
end level_vec_gen;

architecture Behavioral of level_vec_gen is
begin
    process (frame_index, frame_id)
    begin
        -- Update this function to match your requirements
        case frame_index is
            when "000" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0100011100111011010011101100000101011100000110101000111000010000";
                    when "00001" => level_vec_out <= "0100011100111011010011101100100101011100001110101000111000010000";
                    when "00010" => level_vec_out <= "0100011100111011010011101100100101011100001110111000111000010000";
                    when "00011" => level_vec_out <= "0100011100111011010011101100100101011100001110111000111000010000";
                    when "00100" => level_vec_out <= "0101011100111011010011101100100101011100001110111000111000010000";
                    when "00101" => level_vec_out <= "0101011100111011010111101100100101011100001110111000111000010000";
                    when "00110" => level_vec_out <= "0101011100111111010111101100100101011100001110111000111001010001";
                    when "00111" => level_vec_out <= "0101011100111111010111101100100101011100001110111000111001010001";
                    when "01000" => level_vec_out <= "0101011100111111010111101100100101011100001110111000111101110001";
                    when "01001" => level_vec_out <= "0101011100111111010111101100100101111100011110111000111101110001";
                    when "01010" => level_vec_out <= "0101011100111111010111101100100101111100011110111000111101110101";
                    when "01011" => level_vec_out <= "0101011100111111010111101100100101111100011110111001111101110101";
                    when "01100" => level_vec_out <= "0111011100111111010111101110100101111100011110111001111101110101";
                    when "01101" => level_vec_out <= "0111011100111111010111101110100101111100011110111001111101110101";
                    when "01110" => level_vec_out <= "0111011100111111010111101110100101111110011110111001111101110101";
                    when "01111" => level_vec_out <= "0111011100111111010111101110100101111110011110111001111101110101";
                    when "10000" => level_vec_out <= "0111011100111111010111101110100101111110011110111001111101110101";
                    when "10001" => level_vec_out <= "0111011110111111010111101111100101111111011110111001111101110101";
                    when "10010" => level_vec_out <= "1111011110111111010111101111100101111111011111111001111101110101";
                    when "10011" => level_vec_out <= "1111011110111111010111101111100101111111011111111001111101110101";
                    when "10100" => level_vec_out <= "1111011110111111010111101111100101111111011111111001111101110101";
                    when "10101" => level_vec_out <= "1111011110111111010111101111100101111111011111111001111101110101";
                    when "10110" => level_vec_out <= "1111111110111111010111101111100101111111011111111001111101110101";
                    when "10111" => level_vec_out <= "1111111110111111010111101111100101111111011111111001111101110101";
                    when "11000" => level_vec_out <= "1111111110111111010111101111100101111111011111111001111101110101";
                    when "11001" => level_vec_out <= "1111111110111111010111101111100101111111011111111001111101111111";
                    when "11010" => level_vec_out <= "1111111110111111111111101111100101111111011111111001111101111111";
                    when "11011" => level_vec_out <= "1111111110111111111111101111100101111111011111111001111101111111";
                    when "11100" => level_vec_out <= "1111111111111111111111101111100101111111111111111101111101111111";
                    when "11101" => level_vec_out <= "1111111111111111111111101111110101111111111111111101111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111101111111111111111111111111101111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111101111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "001" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1110011110001101101111110101101001101111111011101000110010110010";
                    when "00001" => level_vec_out <= "1110011110001101101111111101101101101111111011101000110010110010";
                    when "00010" => level_vec_out <= "1110011110101101101111111101101101101111111011101000110010110010";
                    when "00011" => level_vec_out <= "1110011110101101101111111101101111101111111011101000110010110010";
                    when "00100" => level_vec_out <= "1110011110101101101111111101101111101111111011101000110010110110";
                    when "00101" => level_vec_out <= "1110011110101101101111111101101111101111111011101000110010110110";
                    when "00110" => level_vec_out <= "1110011110101101101111111101101111101111111011101000110010110110";
                    when "00111" => level_vec_out <= "1110011110101101101111111101101111101111111011101001110010110110";
                    when "01000" => level_vec_out <= "1110011110101101101111111101101111101111111011101001110010110110";
                    when "01001" => level_vec_out <= "1110011110101101101111111101101111101111111011101001110010110110";
                    when "01010" => level_vec_out <= "1110011110101101101111111101101111101111111011101001110010110110";
                    when "01011" => level_vec_out <= "1110011110101101101111111101101111101111111011101001110010110110";
                    when "01100" => level_vec_out <= "1110011110101101101111111101101111101111111011101001110011110110";
                    when "01101" => level_vec_out <= "1110111110101101101111111101101111101111111011101001110011110110";
                    when "01110" => level_vec_out <= "1110111110101101101111111101101111101111111011111001110011110110";
                    when "01111" => level_vec_out <= "1110111110101101101111111101101111101111111011111001110011110110";
                    when "10000" => level_vec_out <= "1110111110101101111111111101101111101111111011111001110011110110";
                    when "10001" => level_vec_out <= "1110111110101101111111111101101111101111111011111001110011110111";
                    when "10010" => level_vec_out <= "1110111110101101111111111101101111101111111011111001110011110111";
                    when "10011" => level_vec_out <= "1110111110101101111111111101101111101111111011111001110011110111";
                    when "10100" => level_vec_out <= "1110111110101101111111111101101111101111111011111001110011110111";
                    when "10101" => level_vec_out <= "1110111110101101111111111101101111101111111011111001110111110111";
                    when "10110" => level_vec_out <= "1110111110101101111111111101101111101111111011111001110111111111";
                    when "10111" => level_vec_out <= "1110111110101111111111111111101111101111111011111001110111111111";
                    when "11000" => level_vec_out <= "1110111110101111111111111111101111101111111011111001110111111111";
                    when "11001" => level_vec_out <= "1110111110101111111111111111101111111111111011111001110111111111";
                    when "11010" => level_vec_out <= "1110111110101111111111111111101111111111111011111001110111111111";
                    when "11011" => level_vec_out <= "1110111110101111111111111111101111111111111111111011110111111111";
                    when "11100" => level_vec_out <= "1110111110101111111111111111101111111111111111111011110111111111";
                    when "11101" => level_vec_out <= "1110111110101111111111111111101111111111111111111011110111111111";
                    when "11110" => level_vec_out <= "1111111110101111111111111111101111111111111111111011110111111111";
                    when "11111" => level_vec_out <= "1111111110101111111111111111111111111111111111111111110111111111";
                when others => null;
                end case;
            when "010" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1100110010101000100100101000110011001011011011000100001111101001";
                    when "00001" => level_vec_out <= "1100110010101000100100101000110011001011011011000100001111101001";
                    when "00010" => level_vec_out <= "1100110010101000100101111001110011001011011011000100001111101001";
                    when "00011" => level_vec_out <= "1100110010101000100101111001110011001011011011000100001111101001";
                    when "00100" => level_vec_out <= "1100110010101000100101111001110011011011011011000100001111101001";
                    when "00101" => level_vec_out <= "1100110010101000100101111001110011011011011011000100001111101101";
                    when "00110" => level_vec_out <= "1100110010101000100101111001110011011011011011000100001111101101";
                    when "00111" => level_vec_out <= "1100110010101001100101111001110011011011011011000100001111101101";
                    when "01000" => level_vec_out <= "1100110010101001100101111001110011011011011011000100011111101101";
                    when "01001" => level_vec_out <= "1100110010101001100101111001110011011011011011000100011111101101";
                    when "01010" => level_vec_out <= "1100110010101011100101111001111011011011111011000100011111101101";
                    when "01011" => level_vec_out <= "1100110010101011100101111001111011011011111011000110011111101101";
                    when "01100" => level_vec_out <= "1100110010101011100101111001111011011011111111000111011111101101";
                    when "01101" => level_vec_out <= "1100110010101011100101111001111011011011111111000111011111101101";
                    when "01110" => level_vec_out <= "1100110010101011100101111001111011011011111111000111011111101101";
                    when "01111" => level_vec_out <= "1110110010101011100101111001111011011011111111000111011111101101";
                    when "10000" => level_vec_out <= "1110110010101011100101111101111011011011111111001111011111101101";
                    when "10001" => level_vec_out <= "1110110010101011100101111101111011011011111111001111011111101101";
                    when "10010" => level_vec_out <= "1110110010101011101101111101111011011011111111011111011111101101";
                    when "10011" => level_vec_out <= "1110110011111011101101111111111011011011111111011111011111101101";
                    when "10100" => level_vec_out <= "1110111011111011101101111111111011011011111111011111011111101101";
                    when "10101" => level_vec_out <= "1110111011111011101111111111111011011011111111011111011111101101";
                    when "10110" => level_vec_out <= "1110111011111011101111111111111011011011111111011111011111101101";
                    when "10111" => level_vec_out <= "1110111011111011101111111111111011111011111111011111011111101101";
                    when "11000" => level_vec_out <= "1110111111111011101111111111111011111011111111011111011111101101";
                    when "11001" => level_vec_out <= "1111111111111011101111111111111011111011111111011111011111101101";
                    when "11010" => level_vec_out <= "1111111111111111101111111111111011111011111111011111011111101111";
                    when "11011" => level_vec_out <= "1111111111111111101111111111111011111011111111011111011111111111";
                    when "11100" => level_vec_out <= "1111111111111111111111111111111011111011111111011111011111111111";
                    when "11101" => level_vec_out <= "1111111111111111111111111111111111111111111111011111011111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111111111011111011111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111011111111111";
                when others => null;
                end case;
            when "011" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0001011001110101101011101010001011101101100111011000100100100011";
                    when "00001" => level_vec_out <= "0001111001110101101011101010001011101101100111011000100100100011";
                    when "00010" => level_vec_out <= "0001111001110101101011101010001011101101100111011000100100100011";
                    when "00011" => level_vec_out <= "0001111001110101101011101010001011101111100111011001100100101011";
                    when "00100" => level_vec_out <= "0001111001110101101011101010001011101111100111011001100100101011";
                    when "00101" => level_vec_out <= "1001111001110101101011101010001011101111100111011001100100101011";
                    when "00110" => level_vec_out <= "1001111001110101101011101010101011101111100111011001100100101011";
                    when "00111" => level_vec_out <= "1001111001110101101111101010101011101111100111011001100100101011";
                    when "01000" => level_vec_out <= "1001111001110101101111101010101011101111100111011101100100101011";
                    when "01001" => level_vec_out <= "1001111001111101101111101110101011101111100111011101100100101011";
                    when "01010" => level_vec_out <= "1011111001111101101111101110101011101111100111011101100100101011";
                    when "01011" => level_vec_out <= "1011111001111101101111101110101111101111100111011101100100101011";
                    when "01100" => level_vec_out <= "1011111001111101101111101110101111101111100111011101100100101011";
                    when "01101" => level_vec_out <= "1011111001111101101111101110101111101111100111011101100101101011";
                    when "01110" => level_vec_out <= "1011111011111101101111101111101111101111101111011101100101101011";
                    when "01111" => level_vec_out <= "1011111111111101101111101111101111101111101111011111101101101011";
                    when "10000" => level_vec_out <= "1011111111111101101111101111101111101111101111111111101101111011";
                    when "10001" => level_vec_out <= "1011111111111101101111101111101111101111101111111111101101111011";
                    when "10010" => level_vec_out <= "1011111111111111101111101111101111101111101111111111101101111011";
                    when "10011" => level_vec_out <= "1011111111111111101111101111111111101111101111111111101101111011";
                    when "10100" => level_vec_out <= "1011111111111111101111101111111111101111101111111111101101111011";
                    when "10101" => level_vec_out <= "1011111111111111101111101111111111101111101111111111101101111011";
                    when "10110" => level_vec_out <= "1011111111111111111111101111111111101111101111111111101101111011";
                    when "10111" => level_vec_out <= "1111111111111111111111101111111111101111101111111111101101111011";
                    when "11000" => level_vec_out <= "1111111111111111111111101111111111101111101111111111101101111011";
                    when "11001" => level_vec_out <= "1111111111111111111111101111111111101111101111111111101101111011";
                    when "11010" => level_vec_out <= "1111111111111111111111101111111111101111101111111111101101111011";
                    when "11011" => level_vec_out <= "1111111111111111111111101111111111101111111111111111101101111011";
                    when "11100" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111101111011";
                    when "11101" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111101111011";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111101111011";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111011";
                when others => null;
                end case;
            when "100" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1100001000101110111101101011110001000011001001111111011010100000";
                    when "00001" => level_vec_out <= "1100001000101110111101101011110001000011001001111111011010100000";
                    when "00010" => level_vec_out <= "1100001000101110111111101011110001000011001001111111011010100000";
                    when "00011" => level_vec_out <= "1100001000101110111111101011110001000011001001111111011010100000";
                    when "00100" => level_vec_out <= "1100001000101110111111101011110011000011001001111111011010100000";
                    when "00101" => level_vec_out <= "1100001000101110111111101011110011000011001001111111011010100000";
                    when "00110" => level_vec_out <= "1100001000101110111111101011110011000011001001111111011010100000";
                    when "00111" => level_vec_out <= "1100001000101110111111101011110011010011001001111111111010100000";
                    when "01000" => level_vec_out <= "1100001000101110111111101011110011010011011001111111111010100000";
                    when "01001" => level_vec_out <= "1100001000111110111111101011110011010011011001111111111010100000";
                    when "01010" => level_vec_out <= "1100001000111110111111101011110011010011011001111111111010100001";
                    when "01011" => level_vec_out <= "1100101000111110111111101011110011110011011001111111111010110001";
                    when "01100" => level_vec_out <= "1100111000111110111111101011110011111011011001111111111010110001";
                    when "01101" => level_vec_out <= "1101111000111110111111101011110011111111011001111111111010110001";
                    when "01110" => level_vec_out <= "1101111000111110111111101011110011111111011001111111111010110001";
                    when "01111" => level_vec_out <= "1101111001111110111111101011110011111111111001111111111010110001";
                    when "10000" => level_vec_out <= "1101111001111110111111101011110011111111111101111111111010110001";
                    when "10001" => level_vec_out <= "1101111001111110111111101011110011111111111101111111111010111001";
                    when "10010" => level_vec_out <= "1101111011111110111111101011110111111111111101111111111010111001";
                    when "10011" => level_vec_out <= "1101111011111110111111101011110111111111111101111111111010111001";
                    when "10100" => level_vec_out <= "1101111011111111111111101011111111111111111101111111111010111001";
                    when "10101" => level_vec_out <= "1101111011111111111111101011111111111111111101111111111010111001";
                    when "10110" => level_vec_out <= "1101111011111111111111101111111111111111111101111111111010111001";
                    when "10111" => level_vec_out <= "1101111011111111111111101111111111111111111101111111111010111001";
                    when "11000" => level_vec_out <= "1101111011111111111111101111111111111111111101111111111011111001";
                    when "11001" => level_vec_out <= "1101111111111111111111101111111111111111111101111111111011111001";
                    when "11010" => level_vec_out <= "1101111111111111111111101111111111111111111111111111111111111001";
                    when "11011" => level_vec_out <= "1101111111111111111111101111111111111111111111111111111111111011";
                    when "11100" => level_vec_out <= "1101111111111111111111111111111111111111111111111111111111111011";
                    when "11101" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "101" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1001001011101010011001100110101010111010011010100000000011101010";
                    when "00001" => level_vec_out <= "1001001011101010011001100110101010111010011010100110000111101010";
                    when "00010" => level_vec_out <= "1001001011101010011001100110101010111010011010100110000111101010";
                    when "00011" => level_vec_out <= "1001001011101010011001100110101010111010011010101110000111101010";
                    when "00100" => level_vec_out <= "1001001011101010011001100110101010111010011010101110000111101110";
                    when "00101" => level_vec_out <= "1001001011101010111001100110101010111011011010101110000111101110";
                    when "00110" => level_vec_out <= "1001001011111010111001100110101010111011011110101110000111101110";
                    when "00111" => level_vec_out <= "1001001011111010111001100110101010111011011110101110000111101110";
                    when "01000" => level_vec_out <= "1001001011111010111001100110101010111011011110101110100111101110";
                    when "01001" => level_vec_out <= "1001001011111010111001100110101010111011011110101110100111101110";
                    when "01010" => level_vec_out <= "1001001011111010111001100110101010111011011110101110100111101110";
                    when "01011" => level_vec_out <= "1101001011111010111001100110101010111011011110101110100111101110";
                    when "01100" => level_vec_out <= "1101001111111010111001100110101010111011011110101110100111101110";
                    when "01101" => level_vec_out <= "1101001111111010111001100111101010111011011110101110100111101110";
                    when "01110" => level_vec_out <= "1101001111111010111001100111101010111011011110101110100111101110";
                    when "01111" => level_vec_out <= "1101001111111011111001100111101010111011011110101110100111101110";
                    when "10000" => level_vec_out <= "1101001111111011111001100111101010111011011110101110100111101110";
                    when "10001" => level_vec_out <= "1101001111111011111001100111101010111011011110101110100111101110";
                    when "10010" => level_vec_out <= "1101001111111011111001100111101010111011011110101110100111101110";
                    when "10011" => level_vec_out <= "1101001111111011111001100111101010111011011110101110100111111110";
                    when "10100" => level_vec_out <= "1101001111111111111001100111101010111011011110101110100111111110";
                    when "10101" => level_vec_out <= "1101001111111111111001100111101010111011011111101111100111111110";
                    when "10110" => level_vec_out <= "1101001111111111111001100111101010111011111111101111100111111110";
                    when "10111" => level_vec_out <= "1101001111111111111001111111101010111011111111101111100111111110";
                    when "11000" => level_vec_out <= "1101101111111111111001111111101010111111111111101111100111111111";
                    when "11001" => level_vec_out <= "1101101111111111111001111111111110111111111111101111100111111111";
                    when "11010" => level_vec_out <= "1101101111111111111011111111111110111111111111101111100111111111";
                    when "11011" => level_vec_out <= "1101101111111111111111111111111110111111111111101111100111111111";
                    when "11100" => level_vec_out <= "1101101111111111111111111111111110111111111111101111100111111111";
                    when "11101" => level_vec_out <= "1101101111111111111111111111111110111111111111101111100111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111110111111111111111111110111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111110111111111";
                when others => null;
                end case;
            when "110" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1010010101000011001011100000110101010111011011100110000111010101";
                    when "00001" => level_vec_out <= "1010010101000011001011100000110101010111011011100110000111010101";
                    when "00010" => level_vec_out <= "1010010101000011001011101000110101010111111011100110000111010101";
                    when "00011" => level_vec_out <= "1010010101000011001011101001110101010111111011100110000111010101";
                    when "00100" => level_vec_out <= "1010010101000111001011101001111101010111111011100110000111010101";
                    when "00101" => level_vec_out <= "1010010101100111001011101001111101010111111011100110001111010101";
                    when "00110" => level_vec_out <= "1010010101100111001011101001111101110111111011100110001111010101";
                    when "00111" => level_vec_out <= "1010010101100111101011101001111101110111111011100110001111010101";
                    when "01000" => level_vec_out <= "1010010101100111101011101101111101110111111011100110011111010101";
                    when "01001" => level_vec_out <= "1010010101100111101011101101111101110111111011100110011111010111";
                    when "01010" => level_vec_out <= "1010010101100111101011101101111101110111111011100110011111010111";
                    when "01011" => level_vec_out <= "1010010111100111101011101101111101110111111011100110011111010111";
                    when "01100" => level_vec_out <= "1010010111100111101011101101111101110111111011100110011111010111";
                    when "01101" => level_vec_out <= "1010010111100111101011101101111101110111111011100110011111110111";
                    when "01110" => level_vec_out <= "1010010111100111101011111101111101110111111011100110011111110111";
                    when "01111" => level_vec_out <= "1010010111100111101011111101111101110111111011100110011111110111";
                    when "10000" => level_vec_out <= "1010010111100111111011111101111101110111111011100110011111110111";
                    when "10001" => level_vec_out <= "1010110111100111111011111101111101110111111011100110011111110111";
                    when "10010" => level_vec_out <= "1010110111100111111011111101111101110111111011101110011111110111";
                    when "10011" => level_vec_out <= "1010110111100111111011111101111101110111111011101110011111111111";
                    when "10100" => level_vec_out <= "1010110111100111111011111101111101110111111111101110011111111111";
                    when "10101" => level_vec_out <= "1011110111100111111011111101111101110111111111101110011111111111";
                    when "10110" => level_vec_out <= "1011110111100111111011111101111101110111111111111111011111111111";
                    when "10111" => level_vec_out <= "1011110111100111111011111101111101111111111111111111111111111111";
                    when "11000" => level_vec_out <= "1011111111100111111011111111111101111111111111111111111111111111";
                    when "11001" => level_vec_out <= "1011111111100111111011111111111101111111111111111111111111111111";
                    when "11010" => level_vec_out <= "1011111111100111111111111111111101111111111111111111111111111111";
                    when "11011" => level_vec_out <= "1111111111101111111111111111111101111111111111111111111111111111";
                    when "11100" => level_vec_out <= "1111111111101111111111111111111101111111111111111111111111111111";
                    when "11101" => level_vec_out <= "1111111111101111111111111111111111111111111111111111111111111111";
                    when "11110" => level_vec_out <= "1111111111101111111111111111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "111" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0101000111001001101111101000000111011010001110100000100001101011";
                    when "00001" => level_vec_out <= "0101000111001001101111101000000111011010001110100000100001101011";
                    when "00010" => level_vec_out <= "0101000111001001101111101000000111011010001110100000100001101011";
                    when "00011" => level_vec_out <= "0101000111001001101111101000100111011011001110100000100001101011";
                    when "00100" => level_vec_out <= "0101000111001001101111101100100111011011001110100000100001101011";
                    when "00101" => level_vec_out <= "0101000111001001101111101100100111011011001110100010100001101011";
                    when "00110" => level_vec_out <= "0101000111011001101111101100100111011011001110100010100001101011";
                    when "00111" => level_vec_out <= "0101010111011001101111101100100111011011001110100010100001101111";
                    when "01000" => level_vec_out <= "0101010111011001101111101100100111011011001110100010100001101111";
                    when "01001" => level_vec_out <= "0101011111011001101111101100100111111011001110100010100001101111";
                    when "01010" => level_vec_out <= "0101011111011001111111101100100111111011001111100010100001101111";
                    when "01011" => level_vec_out <= "0101011111011001111111101100100111111011001111100010100001101111";
                    when "01100" => level_vec_out <= "0101011111011001111111101100100111111011001111100010100001101111";
                    when "01101" => level_vec_out <= "0111011111011001111111111100100111111011001111100010100001101111";
                    when "01110" => level_vec_out <= "1111011111011001111111111100100111111011001111100010101001101111";
                    when "01111" => level_vec_out <= "1111011111011001111111111100100111111011011111100010101001101111";
                    when "10000" => level_vec_out <= "1111011111011001111111111101100111111011011111100010101001101111";
                    when "10001" => level_vec_out <= "1111011111011101111111111101100111111111011111100010101001101111";
                    when "10010" => level_vec_out <= "1111011111011101111111111101100111111111011111100010101001101111";
                    when "10011" => level_vec_out <= "1111011111011101111111111101100111111111011111100010101111101111";
                    when "10100" => level_vec_out <= "1111011111011101111111111101100111111111011111101111101111101111";
                    when "10101" => level_vec_out <= "1111111111011111111111111101100111111111011111101111111111101111";
                    when "10110" => level_vec_out <= "1111111111011111111111111111100111111111011111101111111111101111";
                    when "10111" => level_vec_out <= "1111111111011111111111111111100111111111011111101111111111101111";
                    when "11000" => level_vec_out <= "1111111111011111111111111111100111111111011111101111111111111111";
                    when "11001" => level_vec_out <= "1111111111111111111111111111100111111111011111101111111111111111";
                    when "11010" => level_vec_out <= "1111111111111111111111111111100111111111011111101111111111111111";
                    when "11011" => level_vec_out <= "1111111111111111111111111111100111111111011111101111111111111111";
                    when "11100" => level_vec_out <= "1111111111111111111111111111100111111111011111101111111111111111";
                    when "11101" => level_vec_out <= "1111111111111111111111111111100111111111011111111111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111110111111111011111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111110111111111111111111111111111111111";
                when others => null;
                end case;
            when others => null;
        end case;
    end process;
end Behavioral;