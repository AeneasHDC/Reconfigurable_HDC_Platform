
/**
 * @file class_hvec_gen_hdl.hpp
 * @brief This script generates HDL code for generating high-dimensional class vectors.
 * It is a novel method; for more information, please refer to our paper.
 *
 * @author Saeid Jamili and Marco Angioli
 * @note Author names are listed in alphabetical order.
 * @email <saeid.jamili@uniroma1.it>
 * @email <marco.angioli@uniroma1.it>
 *
 * @contributors
 *
 * @date Created: 24th July 2023
 * @date Last Updated: 23th August 2023
 *
 * @version 1.0.0
 *
 * @institute Sapienza University of Rome
 * @cite https://doi.org/10.xxxx/yyyyy
 *
 * @section DEPENDENCIES
 * - Dependency1: Description or version details.
 * - Dependency2: Description or version details.
 *
 * @section LICENSE
 * This file is part of the Aeneas HyperCompute Platform.
 *
 * Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 *
 * @section CHANGELOG
 * @version 1.0.0-dev - 23th August 2023
 * - Initial release
 *
 * @todo
 * - Complete level vector generator function
 * - Add training
 *
 * @see
 * -
 * -
 * -
 *
 */

module class_hvec_gen #(parameter int DI_PARALLEL_W_BITS = 64) (
  input logic [2:0] frame_id,
  input logic [1:0] frame_index,
  output logic [DI_PARALLEL_W_BITS-1:0] class_vec_out
);
  always_comb begin
    case (frame_id)
      0:
        case (frame_index)
          0:
            class_vec_out = 64'b199971340291990098001991019987199199199058187019919917311619601256419917301779411519712199019601491991141991990531471479590201990199199199199118;
          1:
            class_vec_out = 64'b3611904360021003400361636363601635036363211360241436320331718351336035125362736360022932133053603636363619;
          2:
            class_vec_out = 64'b206507200050019102022020200614020201518190151120160971620520019018201220200101016212042002020202014;
        endcase
      1:
        case (frame_index)
          0:
            class_vec_out = 64'b1991599243199019900901931990019905002300134123019901998383136119019901990028019919919901990018301991996106919991019901991719900;
          1:
            class_vec_out = 64'b363518183603600293536003600001300323203603662021340360360015036363603600350363627025361203603683600;
          2:
            class_vec_out = 64'b2015815200200017152000200100900816020020118713020020002020202002000180202080920502002072000;
        endcase
      2:
        case (frame_index)
          0:
            class_vec_out = 64'b19904151051424199019989240063011500000199199001990000006801210199158199011995901970199680199510419919900196141016501199;
          1:
            class_vec_out = 64'b360302620036236202100501800000363600350000005026036333600366034036603602836360034300310036;
          2:
            class_vec_out = 64'b2002015942012012200801400000202000200000001201702092004201102002080200920200018130180420;
        endcase
      3:
        case (frame_index)
          0:
            class_vec_out = 64'b199147145019918319961621946199001990211140241994818446671681991990017000421991991993111991790199021199199581991990199185069194199396000;
          1:
            class_vec_out = 64'b3672903631365322853600360125020361135122183636003400236363620362903602236362363603619083536155000;
          2:
            class_vec_out = 64'b20790201320181522000200017061931141110142020001600820202030201802002220201202002014111102043000;
        endcase
      4:
        case (frame_index)
          0:
            class_vec_out = 64'b0198195019905919819929836195128167016011219511233199199199981119921741962201995133019274199168199201990581956901580193831970120180291071991080117;
          1:
            class_vec_out = 64'b036310360235360194311331018262681236363647360263680362330312363036003601636301303126330121206263631014;
          2:
            class_vec_out = 64'b0201502001192081071514110131517101120202055200121720200120145201420002006201007014121708705112017017;
        endcase
      5:
        case (frame_index)
          0:
            class_vec_out = 64'b019903201993318917015219919819984701991101991994199148199019901801410199001990943930199199086093801991991991980019919927519819500199116199;
          1:
            class_vec_out = 64'b03605036032333436343672036353636036263603206034036003602830036360180133036363636003636153353400361836;
          2:
            class_vec_out = 64'b02009120620161320172090020152020220720018020150200020017820202001309820202020002020151191900201420;
        endcase
      6:
        case (frame_index)
          0:
            class_vec_out = 64'b584921991590019913199199019919918019919900841991970199121191001111991981919519931991991991991991991997016451193001991990001991311991583199096;
          1:
            class_vec_out = 64'b0189363200363363603636116363600936350362535000036366363603636363636363626355130036360003525363303605;
          2:
            class_vec_out = 64'b2592017002062020020204820200013202002015200070202041920020202020202020819441100202000020122016320013;
        endcase
      7:
        case (frame_index)
          0:
            class_vec_out = 64'b1271024199118199199199199019416199199060419901990199186150199000019915259199199018700761991999612019901990199147199148081991481781981990199199;
          1:
            class_vec_out = 64'b14002363336363636035636360100360360363630360000353433636034005363627503603603623361700363334353603636;
          2:
            class_vec_out = 64'b1000320162020202001442020010220020020111420000017164202001900220209302002002010201302201214172002016;
        endcase
    endcase
  end
endmodule