----
 -- @file level_hvec_gen_hdl.hpp
 -- @brief This script generates HDL code for generating high-dimensional LEVEL vectors.
 -- It is a novel method; for more information, please refer to our paper.
 --
 -- @author Saeid Jamili and Marco Angioli
 -- @note Author names are listed in alphabetical order.
 -- @email <saeid.jamili@uniroma1.it>
 -- @email <marco.angioli@uniroma1.it>
 --
 -- @contributors
 --
 -- @date Created: 24th July 2023
 -- @date Last Updated: 23th August 2023
 --
 -- @version 1.0.0
 --
 -- @institute Sapienza University of Rome
 -- @cite https://doi.org/10.xxxx/yyyyy
 --
 -- @section DEPENDENCIES
 -- - Dependency1: Description or version details.
 -- - Dependency2: Description or version details.
 --
 -- @section LICENSE
 -- This file is part of the Aeneas HyperCompute Platform.
 --
 -- Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 --
 -- @section CHANGELOG
 -- @version 1.0.0-dev - 23th August 2023
 -- - Initial release
 --
 -- @todo
 -- - Complete level vector generator function
 -- - Add training
 --
 -- @see
 -- -
 -- -
 -- -
 --
 --

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity level_vec_gen is
    Port ( level_vec_out : out  STD_LOGIC_VECTOR (63 downto 0);
           frame_index : in  STD_LOGIC_VECTOR (2 downto 0);
           frame_id : in  STD_LOGIC_VECTOR (4 downto 0));
end level_vec_gen;

architecture Behavioral of level_vec_gen is
begin
    process (frame_index, frame_id)
    begin
        -- Update this function to match your requirements
        case frame_index is
            when "000" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0110101101101110010010001111000000100111000011010111000001011111";
                    when "00001" => level_vec_out <= "0110101101101110010010001111000000100111000011010111001001011111";
                    when "00010" => level_vec_out <= "0110101101111110010010011111000010100111000011010111001001011111";
                    when "00011" => level_vec_out <= "0110101101111110010010011111000010100111000011010111001001011111";
                    when "00100" => level_vec_out <= "0110101101111110010010011111000010100111001011010111001001011111";
                    when "00101" => level_vec_out <= "0110101101111110010010011111000010100111101011010111001001011111";
                    when "00110" => level_vec_out <= "0110101101111110010010011111000010100111101011010111001001011111";
                    when "00111" => level_vec_out <= "0110101101111110010110011111000010100111101011010111101001011111";
                    when "01000" => level_vec_out <= "0110101101111110010110011111000010101111101011010111101001011111";
                    when "01001" => level_vec_out <= "0110101101111110010110011111000010101111101011010111101001011111";
                    when "01010" => level_vec_out <= "0110101101111110010110011111000010101111101011010111101001011111";
                    when "01011" => level_vec_out <= "0110101101111110010110011111000010101111101011010111101001111111";
                    when "01100" => level_vec_out <= "0110101101111110010110011111000110101111101011010111101001111111";
                    when "01101" => level_vec_out <= "0110101101111110010110011111000110101111101011010111101001111111";
                    when "01110" => level_vec_out <= "0110101101111110010110011111000110101111101011010111101001111111";
                    when "01111" => level_vec_out <= "0110101101111110010110011111010110101111101011010111101001111111";
                    when "10000" => level_vec_out <= "0110101101111110110110011111010110101111101111010111101001111111";
                    when "10001" => level_vec_out <= "0110101101111110110110011111010110101111101111010111101001111111";
                    when "10010" => level_vec_out <= "0110101101111110110110111111010110101111101111010111101001111111";
                    when "10011" => level_vec_out <= "0110101101111110110110111111010110101111111111010111101001111111";
                    when "10100" => level_vec_out <= "0110101101111110110110111111010110101111111111010111101001111111";
                    when "10101" => level_vec_out <= "0111101101111110110110111111010110101111111111010111101001111111";
                    when "10110" => level_vec_out <= "0111101111111110110110111111010110101111111111011111101001111111";
                    when "10111" => level_vec_out <= "0111101111111110110110111111010110101111111111011111101001111111";
                    when "11000" => level_vec_out <= "0111101111111110110110111111011110101111111111111111101001111111";
                    when "11001" => level_vec_out <= "0111101111111110111110111111011110101111111111111111101001111111";
                    when "11010" => level_vec_out <= "0111101111111110111110111111111110101111111111111111111001111111";
                    when "11011" => level_vec_out <= "0111101111111110111110111111111110101111111111111111111101111111";
                    when "11100" => level_vec_out <= "1111101111111110111110111111111110101111111111111111111101111111";
                    when "11101" => level_vec_out <= "1111111111111110111110111111111111101111111111111111111101111111";
                    when "11110" => level_vec_out <= "1111111111111110111110111111111111101111111111111111111101111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111101111111";
                when others => null;
                end case;
            when "001" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0001110101100101101001011101100100010010001000101000101110010010";
                    when "00001" => level_vec_out <= "0001111101100101101001011101100100010110001000101000101110010010";
                    when "00010" => level_vec_out <= "0001111101100101101001011101100100010110001000101000101110010010";
                    when "00011" => level_vec_out <= "0001111101100101101001011101101100010110001000101000101110010010";
                    when "00100" => level_vec_out <= "1001111101100101101001011101101100010110001010101000101110010010";
                    when "00101" => level_vec_out <= "1001111101100101101001011101101100010110001010101000101110010010";
                    when "00110" => level_vec_out <= "1001111101100101101001011101101100110110001010101100101110010010";
                    when "00111" => level_vec_out <= "1001111101100101101001011101101100110110001010101100101110010010";
                    when "01000" => level_vec_out <= "1001111101101101101101011101101100110110001010101100111110010010";
                    when "01001" => level_vec_out <= "1001111101101101101101011101101101110110101010101100111110010010";
                    when "01010" => level_vec_out <= "1001111101101111101101011101101101110111101010101100111110010011";
                    when "01011" => level_vec_out <= "1101111101101111101101011101101101110111101010101100111110010011";
                    when "01100" => level_vec_out <= "1101111101101111101101011101101101110111111010101100111110010011";
                    when "01101" => level_vec_out <= "1101111101101111101101011101101101110111111110101100111110010011";
                    when "01110" => level_vec_out <= "1101111111101111101101011101101101110111111110101100111110010011";
                    when "01111" => level_vec_out <= "1101111111101111101111011101101101110111111110101100111110010011";
                    when "10000" => level_vec_out <= "1101111111101111101111011101101101110111111110101110111110010011";
                    when "10001" => level_vec_out <= "1101111111101111101111111111101101110111111110111110111110010011";
                    when "10010" => level_vec_out <= "1101111111101111101111111111101111110111111110111110111110010011";
                    when "10011" => level_vec_out <= "1101111111101111101111111111101111110111111110111110111110010011";
                    when "10100" => level_vec_out <= "1101111111101111101111111111101111110111111110111110111110010011";
                    when "10101" => level_vec_out <= "1101111111101111101111111111111111110111111110111110111110010011";
                    when "10110" => level_vec_out <= "1101111111101111101111111111111111110111111110111110111110010011";
                    when "10111" => level_vec_out <= "1101111111101111101111111111111111110111111110111110111110010011";
                    when "11000" => level_vec_out <= "1101111111101111101111111111111111110111111110111110111110110011";
                    when "11001" => level_vec_out <= "1101111111101111101111111111111111110111111110111110111110110011";
                    when "11010" => level_vec_out <= "1111111111101111101111111111111111110111111110111110111110110011";
                    when "11011" => level_vec_out <= "1111111111101111101111111111111111110111111110111110111110110011";
                    when "11100" => level_vec_out <= "1111111111101111101111111111111111110111111110111110111110110111";
                    when "11101" => level_vec_out <= "1111111111101111101111111111111111110111111110111110111110111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111110111111110111111111110111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111110111111111110111111";
                when others => null;
                end case;
            when "010" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0011011100101000010101110001010001011010100101101001110001110111";
                    when "00001" => level_vec_out <= "0011011100101000010101110001010001011010100101101001110001110111";
                    when "00010" => level_vec_out <= "0011011100101000010101110001010001011010100101101001110001110111";
                    when "00011" => level_vec_out <= "0011011100101000010111110001010001011010100101101001110001110111";
                    when "00100" => level_vec_out <= "0011011100101000010111110001010001011010100101101001110001110111";
                    when "00101" => level_vec_out <= "0011011100111000010111110001010001011010110101101001110001110111";
                    when "00110" => level_vec_out <= "0011011100111000010111110001010001011010110101101001110001110111";
                    when "00111" => level_vec_out <= "0011011100111000010111110001010001011010110101101001110001110111";
                    when "01000" => level_vec_out <= "0011011100111000010111110001010001011010110101101001110101110111";
                    when "01001" => level_vec_out <= "0111011100111000010111110001010001011010110101101001110101110111";
                    when "01010" => level_vec_out <= "0111011100111000010111111001010001011010110101101001110101110111";
                    when "01011" => level_vec_out <= "0111011100111000010111111001010001011010110101101011110101110111";
                    when "01100" => level_vec_out <= "0111011100111000010111111001010001011010110101101011110101110111";
                    when "01101" => level_vec_out <= "0111011100111000010111111001010101111010110101101011110101110111";
                    when "01110" => level_vec_out <= "0111011100111000010111111001010101111010110111101011110101110111";
                    when "01111" => level_vec_out <= "0111011100111000010111111001010101111010110111101011110101110111";
                    when "10000" => level_vec_out <= "0111011100111010010111111001010101111010110111101011110101110111";
                    when "10001" => level_vec_out <= "0111011110111010010111111001010101111010110111101011110101110111";
                    when "10010" => level_vec_out <= "0111011110111010010111111001010101111010110111111011110101110111";
                    when "10011" => level_vec_out <= "1111011110111110010111111001110101111010110111111011110101110111";
                    when "10100" => level_vec_out <= "1111011110111110011111111001110101111010110111111111111111111111";
                    when "10101" => level_vec_out <= "1111011110111110011111111001110101111110110111111111111111111111";
                    when "10110" => level_vec_out <= "1111011110111111011111111001110101111110111111111111111111111111";
                    when "10111" => level_vec_out <= "1111011110111111011111111001111101111110111111111111111111111111";
                    when "11000" => level_vec_out <= "1111111110111111011111111001111101111110111111111111111111111111";
                    when "11001" => level_vec_out <= "1111111110111111011111111001111101111110111111111111111111111111";
                    when "11010" => level_vec_out <= "1111111110111111011111111001111101111110111111111111111111111111";
                    when "11011" => level_vec_out <= "1111111110111111011111111001111101111110111111111111111111111111";
                    when "11100" => level_vec_out <= "1111111110111111011111111011111101111110111111111111111111111111";
                    when "11101" => level_vec_out <= "1111111110111111011111111011111101111111111111111111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111011111111011111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "011" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0101000101100100000100111011101110011011100100101110011010111100";
                    when "00001" => level_vec_out <= "0101000101100100000100111011101110011011100100101110011010111100";
                    when "00010" => level_vec_out <= "0101000101100100000100111011101110011011101100101110011010111100";
                    when "00011" => level_vec_out <= "0101000101100100000100111011101110011011101100101111011010111100";
                    when "00100" => level_vec_out <= "0101000101100100010100111011101110011011101100101111011010111100";
                    when "00101" => level_vec_out <= "0101001101100100010100111011101110011011101100101111011010111100";
                    when "00110" => level_vec_out <= "0111001101100100010100111011101110011011101100101111011010111100";
                    when "00111" => level_vec_out <= "0111001101100100010100111011101110011011101100101111011010111100";
                    when "01000" => level_vec_out <= "0111001101100100010100111011101110011011101100101111011010111100";
                    when "01001" => level_vec_out <= "0111001101100100010100111011101110011011101100101111011010111100";
                    when "01010" => level_vec_out <= "0111001101100101010100111011101110011011101100101111011010111100";
                    when "01011" => level_vec_out <= "0111001101100101010101111111101110011011101100101111011010111100";
                    when "01100" => level_vec_out <= "0111001101100101010101111111111110011011101100101111011010111100";
                    when "01101" => level_vec_out <= "0111001101100101010101111111111110011011101100101111011010111100";
                    when "01110" => level_vec_out <= "0111001101100101010101111111111110011011101110101111011010111100";
                    when "01111" => level_vec_out <= "0111001101100101010101111111111110011011111110101111011010111101";
                    when "10000" => level_vec_out <= "0111001101100101010101111111111110011011111110101111011010111101";
                    when "10001" => level_vec_out <= "0111001101100101010111111111111110011011111110101111011010111101";
                    when "10010" => level_vec_out <= "0111101101100101010111111111111110111011111110101111011010111101";
                    when "10011" => level_vec_out <= "0111101101100101010111111111111110111011111110101111011010111111";
                    when "10100" => level_vec_out <= "0111101101100101010111111111111110111011111110101111011010111111";
                    when "10101" => level_vec_out <= "0111101111100101011111111111111110111011111110101111011010111111";
                    when "10110" => level_vec_out <= "0111101111100101011111111111111110111011111110101111011010111111";
                    when "10111" => level_vec_out <= "0111101111100101111111111111111110111011111110111111011010111111";
                    when "11000" => level_vec_out <= "0111101111101101111111111111111110111011111110111111011010111111";
                    when "11001" => level_vec_out <= "0111101111101111111111111111111110111111111110111111011011111111";
                    when "11010" => level_vec_out <= "0111101111101111111111111111111110111111111110111111011111111111";
                    when "11011" => level_vec_out <= "1111101111101111111111111111111110111111111111111111011111111111";
                    when "11100" => level_vec_out <= "1111101111101111111111111111111110111111111111111111011111111111";
                    when "11101" => level_vec_out <= "1111101111101111111111111111111110111111111111111111111111111111";
                    when "11110" => level_vec_out <= "1111101111101111111111111111111110111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111101111101111111111111111111110111111111111111111111111111111";
                when others => null;
                end case;
            when "100" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0111000010101010011111110011010001110100110000100111101011100010";
                    when "00001" => level_vec_out <= "1111001010101010011111110011010001110100110000100111101011100010";
                    when "00010" => level_vec_out <= "1111001010101010011111110011010001110100110010100111101011100010";
                    when "00011" => level_vec_out <= "1111001010111010011111110011010001110100110010100111111011100010";
                    when "00100" => level_vec_out <= "1111001010111011011111110011010001110100110010101111111011100010";
                    when "00101" => level_vec_out <= "1111001010111011011111110011010001110100110010101111111011100010";
                    when "00110" => level_vec_out <= "1111001010111011011111110011010001110100111011101111111011100010";
                    when "00111" => level_vec_out <= "1111001010111011011111110111010001110100111011101111111011101010";
                    when "01000" => level_vec_out <= "1111001010111011011111110111010001110100111011101111111011101010";
                    when "01001" => level_vec_out <= "1111001010111011011111110111010001110101111011101111111011101010";
                    when "01010" => level_vec_out <= "1111101010111011011111110111010001110101111011101111111011101010";
                    when "01011" => level_vec_out <= "1111101010111011011111110111010001110101111011101111111011101010";
                    when "01100" => level_vec_out <= "1111101010111011011111110111010101110101111111101111111011101010";
                    when "01101" => level_vec_out <= "1111101010111011011111110111010101110101111111101111111011101010";
                    when "01110" => level_vec_out <= "1111101010111011011111110111110101110101111111101111111011101010";
                    when "01111" => level_vec_out <= "1111101010111011011111110111111101110101111111101111111011101010";
                    when "10000" => level_vec_out <= "1111101010111011011111110111111101110101111111101111111011101010";
                    when "10001" => level_vec_out <= "1111101010111011011111110111111101110101111111101111111011101010";
                    when "10010" => level_vec_out <= "1111101010111011011111110111111101110101111111101111111011101010";
                    when "10011" => level_vec_out <= "1111101010111011011111110111111101110101111111101111111011101010";
                    when "10100" => level_vec_out <= "1111101010111111011111110111111101110101111111101111111011101010";
                    when "10101" => level_vec_out <= "1111101010111111011111110111111101110101111111101111111011101010";
                    when "10110" => level_vec_out <= "1111101010111111011111111111111101111101111111101111111011101010";
                    when "10111" => level_vec_out <= "1111101010111111011111111111111101111101111111101111111111101010";
                    when "11000" => level_vec_out <= "1111101011111111011111111111111101111111111111101111111111101010";
                    when "11001" => level_vec_out <= "1111101011111111011111111111111101111111111111101111111111101011";
                    when "11010" => level_vec_out <= "1111111011111111111111111111111101111111111111101111111111101011";
                    when "11011" => level_vec_out <= "1111111011111111111111111111111101111111111111101111111111101011";
                    when "11100" => level_vec_out <= "1111111111111111111111111111111101111111111111101111111111101111";
                    when "11101" => level_vec_out <= "1111111111111111111111111111111111111111111111101111111111101111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111111111101111111111101111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "101" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0010101110000101000110110100010001010101000011001001100011010101";
                    when "00001" => level_vec_out <= "0010101110000101000110110100010001011101000011001001100011010101";
                    when "00010" => level_vec_out <= "0010101110000101000110110100010001011101000011001011100011010101";
                    when "00011" => level_vec_out <= "0010101110100101000110110100010001011101000011001011100011010101";
                    when "00100" => level_vec_out <= "0010101110100101000110110100010001011101000011001011100011010101";
                    when "00101" => level_vec_out <= "0010101110100101000110110100010001011101000011001011100011010101";
                    when "00110" => level_vec_out <= "1010101110100101000110110110010001011101000011001011100011010101";
                    when "00111" => level_vec_out <= "1010101110100101000110110110010001011101000011001011100011010101";
                    when "01000" => level_vec_out <= "1010101110110101000110110110010001011101000011001011100011010101";
                    when "01001" => level_vec_out <= "1010101110110101000110110110010001011101000011001111100011110101";
                    when "01010" => level_vec_out <= "1010101110110101000110110110111001011101000011001111100011110101";
                    when "01011" => level_vec_out <= "1010101110110101000110110110111001111101000011001111100011110101";
                    when "01100" => level_vec_out <= "1010101110110101000110111110111001111101000011001111100011110101";
                    when "01101" => level_vec_out <= "1010101110110101000110111110111101111101001011001111100011110101";
                    when "01110" => level_vec_out <= "1010101110110101000110111110111101111101001011001111100011110101";
                    when "01111" => level_vec_out <= "1010101110110101000110111110111101111101001011101111100011110101";
                    when "10000" => level_vec_out <= "1010101110110101000110111110111101111111001011101111100111110101";
                    when "10001" => level_vec_out <= "1010101110110101000110111110111101111111011011101111100111110101";
                    when "10010" => level_vec_out <= "1010101110110101001110111110111101111111011011101111110111110101";
                    when "10011" => level_vec_out <= "1010101110110101001111111111111101111111011011101111110111110101";
                    when "10100" => level_vec_out <= "1010101110110101001111111111111101111111011011101111110111110101";
                    when "10101" => level_vec_out <= "1010101110110101001111111111111101111111011011101111110111111101";
                    when "10110" => level_vec_out <= "1010101110110101001111111111111101111111011011101111110111111101";
                    when "10111" => level_vec_out <= "1011111110110101001111111111111101111111011011101111110111111101";
                    when "11000" => level_vec_out <= "1011111110110101001111111111111101111111011011101111110111111101";
                    when "11001" => level_vec_out <= "1011111111110101001111111111111101111111011011101111110111111101";
                    when "11010" => level_vec_out <= "1011111111110101001111111111111111111111011011101111110111111101";
                    when "11011" => level_vec_out <= "1011111111110101001111111111111111111111011111101111111111111111";
                    when "11100" => level_vec_out <= "1011111111111101001111111111111111111111111111101111111111111111";
                    when "11101" => level_vec_out <= "1111111111111101001111111111111111111111111111101111111111111111";
                    when "11110" => level_vec_out <= "1111111111111101011111111111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111101011111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "110" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1001001011101000010111101100100110110100011100000001101001001010";
                    when "00001" => level_vec_out <= "1001001011101000010111111100100110110101011100000001101001001010";
                    when "00010" => level_vec_out <= "1001001011101000010111111100110110110101011100000001101001001010";
                    when "00011" => level_vec_out <= "1001001011101000010111111100110110110101011100000001101001001010";
                    when "00100" => level_vec_out <= "1001001011111000010111111100110110110101011100000001101001001010";
                    when "00101" => level_vec_out <= "1001101011111000010111111111110110110101011100000001101001001010";
                    when "00110" => level_vec_out <= "1001101011111000010111111111110110110111011100000001101001001010";
                    when "00111" => level_vec_out <= "1001101111111000010111111111110110110111111100000001101001001010";
                    when "01000" => level_vec_out <= "1001101111111000011111111111110110110111111101000001101001001010";
                    when "01001" => level_vec_out <= "1001101111111000011111111111110110110111111101000001101001001010";
                    when "01010" => level_vec_out <= "1001101111111000011111111111110110110111111101000001101001001010";
                    when "01011" => level_vec_out <= "1001101111111010011111111111110110110111111101000101101001001010";
                    when "01100" => level_vec_out <= "1001101111111010011111111111110110110111111101000101101001101010";
                    when "01101" => level_vec_out <= "1011101111111110011111111111110110110111111101010101101001101010";
                    when "01110" => level_vec_out <= "1011101111111110111111111111110110110111111101010101101001101010";
                    when "01111" => level_vec_out <= "1011111111111110111111111111110110110111111101010101101001111010";
                    when "10000" => level_vec_out <= "1011111111111111111111111111110110110111111101010101101001111010";
                    when "10001" => level_vec_out <= "1011111111111111111111111111110110110111111101110101101001111010";
                    when "10010" => level_vec_out <= "1011111111111111111111111111110110110111111101110101101001111010";
                    when "10011" => level_vec_out <= "1011111111111111111111111111110110110111111101110101101101111010";
                    when "10100" => level_vec_out <= "1111111111111111111111111111110110110111111101110101101111111010";
                    when "10101" => level_vec_out <= "1111111111111111111111111111110110110111111101110101111111111010";
                    when "10110" => level_vec_out <= "1111111111111111111111111111110110110111111101110111111111111110";
                    when "10111" => level_vec_out <= "1111111111111111111111111111110110111111111111110111111111111110";
                    when "11000" => level_vec_out <= "1111111111111111111111111111110110111111111111110111111111111110";
                    when "11001" => level_vec_out <= "1111111111111111111111111111110110111111111111110111111111111110";
                    when "11010" => level_vec_out <= "1111111111111111111111111111110110111111111111110111111111111110";
                    when "11011" => level_vec_out <= "1111111111111111111111111111110110111111111111110111111111111111";
                    when "11100" => level_vec_out <= "1111111111111111111111111111111110111111111111110111111111111111";
                    when "11101" => level_vec_out <= "1111111111111111111111111111111111111111111111110111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "111" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1111100110110111011110001010101110111101101011011010110110001111";
                    when "00001" => level_vec_out <= "1111100110110111011110001010101110111101101011011010110110001111";
                    when "00010" => level_vec_out <= "1111100110110111011110001010101110111101101011011110110110001111";
                    when "00011" => level_vec_out <= "1111101110110111011111001010101110111101101011011110110110001111";
                    when "00100" => level_vec_out <= "1111101110110111011111001010101110111101101011011111110110001111";
                    when "00101" => level_vec_out <= "1111101110110111011111001010101111111101101011011111110110001111";
                    when "00110" => level_vec_out <= "1111101110110111011111001010101111111101101011011111110110001111";
                    when "00111" => level_vec_out <= "1111101110110111011111001010101111111101101111111111110110001111";
                    when "01000" => level_vec_out <= "1111101110110111011111001010101111111101101111111111110110001111";
                    when "01001" => level_vec_out <= "1111111110110111111111001010101111111101101111111111110110001111";
                    when "01010" => level_vec_out <= "1111111110110111111111001010101111111101101111111111110110001111";
                    when "01011" => level_vec_out <= "1111111110110111111111001010101111111101101111111111110110001111";
                    when "01100" => level_vec_out <= "1111111110110111111111001011101111111101101111111111110110001111";
                    when "01101" => level_vec_out <= "1111111110110111111111001011101111111101101111111111110110001111";
                    when "01110" => level_vec_out <= "1111111110110111111111001011101111111111101111111111110111011111";
                    when "01111" => level_vec_out <= "1111111110110111111111001011101111111111101111111111110111011111";
                    when "10000" => level_vec_out <= "1111111110110111111111101011101111111111101111111111110111011111";
                    when "10001" => level_vec_out <= "1111111110110111111111111011101111111111101111111111110111011111";
                    when "10010" => level_vec_out <= "1111111110110111111111111011101111111111101111111111111111011111";
                    when "10011" => level_vec_out <= "1111111110110111111111111011101111111111101111111111111111011111";
                    when "10100" => level_vec_out <= "1111111110110111111111111011101111111111101111111111111111011111";
                    when "10101" => level_vec_out <= "1111111110110111111111111011101111111111101111111111111111111111";
                    when "10110" => level_vec_out <= "1111111110110111111111111011101111111111101111111111111111111111";
                    when "10111" => level_vec_out <= "1111111110110111111111111011101111111111101111111111111111111111";
                    when "11000" => level_vec_out <= "1111111110110111111111111111101111111111101111111111111111111111";
                    when "11001" => level_vec_out <= "1111111111111111111111111111101111111111101111111111111111111111";
                    when "11010" => level_vec_out <= "1111111111111111111111111111101111111111111111111111111111111111";
                    when "11011" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "11100" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "11101" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when others => null;
        end case;
    end process;
end Behavioral;