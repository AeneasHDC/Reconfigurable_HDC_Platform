----
 -- @file level_hvec_gen_hdl.hpp
 -- @brief This script generates HDL code for generating high-dimensional LEVEL vectors.
 -- It is a novel method; for more information, please refer to our paper.
 --
 -- @author Saeid Jamili and Marco Angioli
 -- @note Author names are listed in alphabetical order.
 -- @email <saeid.jamili@uniroma1.it>
 -- @email <marco.angioli@uniroma1.it>
 --
 -- @contributors
 --
 -- @date Created: 24th July 2023
 -- @date Last Updated: 23th August 2023
 --
 -- @version 1.0.0
 --
 -- @institute Sapienza University of Rome
 -- @cite https://doi.org/10.xxxx/yyyyy
 --
 -- @section DEPENDENCIES
 -- - Dependency1: Description or version details.
 -- - Dependency2: Description or version details.
 --
 -- @section LICENSE
 -- This file is part of the Aeneas HyperCompute Platform.
 --
 -- Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 --
 -- @section CHANGELOG
 -- @version 1.0.0-dev - 23th August 2023
 -- - Initial release
 --
 -- @todo
 -- - Complete level vector generator function
 -- - Add training
 --
 -- @see
 -- -
 -- -
 -- -
 --
 --

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity level_vec_gen is
    Port ( level_vec_out : out  STD_LOGIC_VECTOR (63 downto 0);
           frame_index : in  STD_LOGIC_VECTOR (2 downto 0);
           frame_id : in  STD_LOGIC_VECTOR (4 downto 0));
end level_vec_gen;

architecture Behavioral of level_vec_gen is
begin
    process (frame_index, frame_id)
    begin
        -- Update this function to match your requirements
        case frame_index is
            when "000" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1110000000001001111110100000001000001011111110001010101010101100";
                    when "00001" => level_vec_out <= "1110000000001001111110100000001000001011111111001010101010101100";
                    when "00010" => level_vec_out <= "1110000000001001111110100000001000001011111111001010101010101100";
                    when "00011" => level_vec_out <= "1110000000001001111110100000001010001011111111001010111010101100";
                    when "00100" => level_vec_out <= "1110000000001001111110100000001010001011111111101010111010101100";
                    when "00101" => level_vec_out <= "1110000000001001111110100000001010001011111111101010111010101100";
                    when "00110" => level_vec_out <= "1110000100001001111110100000001010001011111111111010111010101100";
                    when "00111" => level_vec_out <= "1110000100001001111110100000001010001011111111111010111010101100";
                    when "01000" => level_vec_out <= "1111000100001001111110100000001010001011111111111110111010101100";
                    when "01001" => level_vec_out <= "1111000100001101111110100000001010001011111111111110111010101100";
                    when "01010" => level_vec_out <= "1111000100001101111110100000001010001011111111111110111010111100";
                    when "01011" => level_vec_out <= "1111000100101101111110100000001010001011111111111110111010111101";
                    when "01100" => level_vec_out <= "1111000100101101111111110000001010001011111111111110111010111101";
                    when "01101" => level_vec_out <= "1111000100101101111111110000001010001011111111111111111010111101";
                    when "01110" => level_vec_out <= "1111000100101101111111110000001010001011111111111111111010111101";
                    when "01111" => level_vec_out <= "1111000100101101111111110000001010001011111111111111111010111101";
                    when "10000" => level_vec_out <= "1111100100101101111111111000001010001011111111111111111110111101";
                    when "10001" => level_vec_out <= "1111100100101101111111111000001010101011111111111111111110111101";
                    when "10010" => level_vec_out <= "1111100100101101111111111000011010101011111111111111111110111111";
                    when "10011" => level_vec_out <= "1111101100101111111111111000011010101111111111111111111110111111";
                    when "10100" => level_vec_out <= "1111101100101111111111111001011010101111111111111111111110111111";
                    when "10101" => level_vec_out <= "1111101100101111111111111001111010101111111111111111111111111111";
                    when "10110" => level_vec_out <= "1111101100101111111111111001111011101111111111111111111111111111";
                    when "10111" => level_vec_out <= "1111101100101111111111111101111011101111111111111111111111111111";
                    when "11000" => level_vec_out <= "1111101100101111111111111101111011101111111111111111111111111111";
                    when "11001" => level_vec_out <= "1111101100101111111111111101111111101111111111111111111111111111";
                    when "11010" => level_vec_out <= "1111111100101111111111111111111111101111111111111111111111111111";
                    when "11011" => level_vec_out <= "1111111100101111111111111111111111101111111111111111111111111111";
                    when "11100" => level_vec_out <= "1111111100101111111111111111111111101111111111111111111111111111";
                    when "11101" => level_vec_out <= "1111111100101111111111111111111111101111111111111111111111111111";
                    when "11110" => level_vec_out <= "1111111110111111111111111111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111110111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "001" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1001111011001110000101100000010000101110100001010101011010000001";
                    when "00001" => level_vec_out <= "1001111011001110000101100000010000101110100001010101011010000001";
                    when "00010" => level_vec_out <= "1001111011001110001101100000010000101110100001010101011011000001";
                    when "00011" => level_vec_out <= "1001111011001110001101100000010000101110100001010101111011000001";
                    when "00100" => level_vec_out <= "1001111011001110001101100000010000101110100001010101111011000001";
                    when "00101" => level_vec_out <= "1001111011001110001101100000010000101110100001010101111011000001";
                    when "00110" => level_vec_out <= "1001111011001110001101100010010000101110100001011101111011100001";
                    when "00111" => level_vec_out <= "1101111011001110001101100010010010101110100001011101111011100001";
                    when "01000" => level_vec_out <= "1101111011001110001101100010010010101110100001011101111011100001";
                    when "01001" => level_vec_out <= "1101111011001110101101100110010010101110100001011101111011100001";
                    when "01010" => level_vec_out <= "1101111011001110101111100110010010101110100001011101111011100001";
                    when "01011" => level_vec_out <= "1101111011001110101111100111010010101110100001011101111011100001";
                    when "01100" => level_vec_out <= "1101111011001110101111110111011010101110100001011101111011100001";
                    when "01101" => level_vec_out <= "1101111011001110101111110111011010101110100011011101111011100001";
                    when "01110" => level_vec_out <= "1101111011001110101111110111111010101110100011011101111011100001";
                    when "01111" => level_vec_out <= "1101111011001110111111110111111010101110110011011101111011100001";
                    when "10000" => level_vec_out <= "1101111011001110111111110111111010101110110011111101111011100001";
                    when "10001" => level_vec_out <= "1101111011001110111111110111111010101110111011111101111011100001";
                    when "10010" => level_vec_out <= "1101111011011110111111110111111010101110111011111101111111100001";
                    when "10011" => level_vec_out <= "1101111011011110111111110111111010111110111011111101111111100001";
                    when "10100" => level_vec_out <= "1101111011011110111111110111111010111110111011111101111111100001";
                    when "10101" => level_vec_out <= "1101111011011110111111110111111010111110111111111101111111100001";
                    when "10110" => level_vec_out <= "1101111011011110111111111111111010111110111111111101111111100101";
                    when "10111" => level_vec_out <= "1111111011011110111111111111111011111110111111111101111111100101";
                    when "11000" => level_vec_out <= "1111111011011110111111111111111011111111111111111101111111100101";
                    when "11001" => level_vec_out <= "1111111011011111111111111111111011111111111111111101111111100111";
                    when "11010" => level_vec_out <= "1111111011011111111111111111111011111111111111111101111111110111";
                    when "11011" => level_vec_out <= "1111111111011111111111111111111011111111111111111101111111110111";
                    when "11100" => level_vec_out <= "1111111111111111111111111111111111111111111111111101111111110111";
                    when "11101" => level_vec_out <= "1111111111111111111111111111111111111111111111111101111111110111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111111111111101111111110111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111110111";
                when others => null;
                end case;
            when "010" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1010011000011111110011011111100011001010110111101011001011000000";
                    when "00001" => level_vec_out <= "1010011000011111110011011111100011001010110111101011001011000000";
                    when "00010" => level_vec_out <= "1010011000011111110011011111100011001010111111101011001011000000";
                    when "00011" => level_vec_out <= "1010011000011111110011011111100011001010111111101011001011000000";
                    when "00100" => level_vec_out <= "1010011000011111110011011111100011001010111111101011001011000000";
                    when "00101" => level_vec_out <= "1010011000011111110011011111100011001010111111101011001111000000";
                    when "00110" => level_vec_out <= "1010011000011111110011011111100011001010111111111011001111001000";
                    when "00111" => level_vec_out <= "1010011000011111110011011111100011001010111111111011001111001010";
                    when "01000" => level_vec_out <= "1011011000011111110011111111100011001010111111111111001111001010";
                    when "01001" => level_vec_out <= "1011011000011111110011111111100011001010111111111111001111001010";
                    when "01010" => level_vec_out <= "1011011000011111110011111111100011001010111111111111001111001010";
                    when "01011" => level_vec_out <= "1011011000011111111011111111100011001010111111111111001111001010";
                    when "01100" => level_vec_out <= "1011111000011111111011111111100011001110111111111111001111001010";
                    when "01101" => level_vec_out <= "1011111000011111111011111111100011001110111111111111001111001010";
                    when "01110" => level_vec_out <= "1011111000011111111011111111100011011110111111111111001111001010";
                    when "01111" => level_vec_out <= "1011111000111111111111111111100011011110111111111111001111001010";
                    when "10000" => level_vec_out <= "1011111100111111111111111111100011011110111111111111001111001010";
                    when "10001" => level_vec_out <= "1011111100111111111111111111100011011110111111111111001111001010";
                    when "10010" => level_vec_out <= "1011111100111111111111111111100011011110111111111111001111001010";
                    when "10011" => level_vec_out <= "1011111101111111111111111111100111011110111111111111001111001010";
                    when "10100" => level_vec_out <= "1011111101111111111111111111110111011110111111111111011111001010";
                    when "10101" => level_vec_out <= "1111111111111111111111111111110111011110111111111111011111001010";
                    when "10110" => level_vec_out <= "1111111111111111111111111111110111111110111111111111011111101010";
                    when "10111" => level_vec_out <= "1111111111111111111111111111110111111110111111111111011111101110";
                    when "11000" => level_vec_out <= "1111111111111111111111111111111111111110111111111111011111101110";
                    when "11001" => level_vec_out <= "1111111111111111111111111111111111111110111111111111011111101110";
                    when "11010" => level_vec_out <= "1111111111111111111111111111111111111110111111111111011111101110";
                    when "11011" => level_vec_out <= "1111111111111111111111111111111111111111111111111111011111111110";
                    when "11100" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111110";
                    when "11101" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111110";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111110";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111110";
                when others => null;
                end case;
            when "011" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0011010011100110000001011101111111100011011011100001110111111000";
                    when "00001" => level_vec_out <= "0011010011100110000001011101111111100011011111100001110111111000";
                    when "00010" => level_vec_out <= "0011010011100110001001011101111111100011011111100001110111111000";
                    when "00011" => level_vec_out <= "0011010011101110001001011101111111100011011111100001110111111000";
                    when "00100" => level_vec_out <= "0011010011101110001001011101111111100011011111100001110111111000";
                    when "00101" => level_vec_out <= "0011010011101110001001011101111111110011011111100011110111111000";
                    when "00110" => level_vec_out <= "0011010011101110001001011101111111110011011111100011110111111000";
                    when "00111" => level_vec_out <= "0011010011101110001001011101111111110111011111100011110111111000";
                    when "01000" => level_vec_out <= "0011010011101110001001011101111111110111011111100011110111111000";
                    when "01001" => level_vec_out <= "0011010011101110001001011101111111111111011111100011110111111000";
                    when "01010" => level_vec_out <= "0011010011101110001001011101111111111111011111100011110111111001";
                    when "01011" => level_vec_out <= "0011011011101110001001011101111111111111011111100011110111111001";
                    when "01100" => level_vec_out <= "0011011011101110001001011101111111111111011111100011110111111011";
                    when "01101" => level_vec_out <= "0011011011101110001001011101111111111111011111100011110111111011";
                    when "01110" => level_vec_out <= "0011011011101110011001011101111111111111011111100011110111111011";
                    when "01111" => level_vec_out <= "0011011011101111011001011101111111111111011111100011110111111011";
                    when "10000" => level_vec_out <= "0011111011101111011001011101111111111111011111100011110111111011";
                    when "10001" => level_vec_out <= "0011111011101111011001011101111111111111111111101011110111111011";
                    when "10010" => level_vec_out <= "0011111011101111011001011111111111111111111111101011110111111011";
                    when "10011" => level_vec_out <= "0011111011101111011001011111111111111111111111101011110111111011";
                    when "10100" => level_vec_out <= "0111111011101111011001011111111111111111111111101011110111111011";
                    when "10101" => level_vec_out <= "0111111011101111011001011111111111111111111111101011110111111011";
                    when "10110" => level_vec_out <= "0111111011101111011001011111111111111111111111101011110111111011";
                    when "10111" => level_vec_out <= "0111111011101111011001011111111111111111111111101011110111111011";
                    when "11000" => level_vec_out <= "0111111011101111011001011111111111111111111111101011110111111011";
                    when "11001" => level_vec_out <= "0111111011101111011001011111111111111111111111101011110111111011";
                    when "11010" => level_vec_out <= "0111111011101111011101011111111111111111111111101011110111111011";
                    when "11011" => level_vec_out <= "0111111011101111011111011111111111111111111111101011110111111111";
                    when "11100" => level_vec_out <= "0111111011111111011111011111111111111111111111101011110111111111";
                    when "11101" => level_vec_out <= "1111111011111111011111111111111111111111111111101011111111111111";
                    when "11110" => level_vec_out <= "1111111111111111011111111111111111111111111111101111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111101111111111111111";
                when others => null;
                end case;
            when "100" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1100010101100100110101010000010101000111111110100011100001011110";
                    when "00001" => level_vec_out <= "1100010101100100110101110000010101000111111110100011100001011110";
                    when "00010" => level_vec_out <= "1110010101100100110101110000010101000111111111100011100001011110";
                    when "00011" => level_vec_out <= "1110010101100110110101110000010101000111111111100011100001011110";
                    when "00100" => level_vec_out <= "1110010101101110110101110000010111000111111111100111100001011110";
                    when "00101" => level_vec_out <= "1110010101101110110101110000010111000111111111100111100001011110";
                    when "00110" => level_vec_out <= "1110010101101110110101110000010111000111111111100111100001011110";
                    when "00111" => level_vec_out <= "1110010101101110110101110000010111000111111111100111101001011110";
                    when "01000" => level_vec_out <= "1110010101101110110101110000110111000111111111100111101001011110";
                    when "01001" => level_vec_out <= "1110010101101110110101110001110111000111111111100111101001011110";
                    when "01010" => level_vec_out <= "1110010101101110110101110001110111010111111111100111101001011110";
                    when "01011" => level_vec_out <= "1110010101101110110101110001110111010111111111100111101001011110";
                    when "01100" => level_vec_out <= "1110010101101110110101110001110111010111111111100111101001011110";
                    when "01101" => level_vec_out <= "1110010101101110110101110001110111010111111111100111101001011110";
                    when "01110" => level_vec_out <= "1110010101101110110101110001110111010111111111100111101001011111";
                    when "01111" => level_vec_out <= "1110010101101110110111110001110111010111111111101111101001011111";
                    when "10000" => level_vec_out <= "1110110101101110110111110001110111010111111111101111101001011111";
                    when "10001" => level_vec_out <= "1110110101101111110111110001110111010111111111101111101001111111";
                    when "10010" => level_vec_out <= "1110110101101111110111110001110111010111111111101111101001111111";
                    when "10011" => level_vec_out <= "1110110101101111110111110001110111010111111111101111101001111111";
                    when "10100" => level_vec_out <= "1110110101101111110111110001110111010111111111101111111001111111";
                    when "10101" => level_vec_out <= "1110110111101111110111110001110111010111111111101111111001111111";
                    when "10110" => level_vec_out <= "1110110111101111110111110001110111110111111111101111111001111111";
                    when "10111" => level_vec_out <= "1111110111101111110111110001110111110111111111101111111001111111";
                    when "11000" => level_vec_out <= "1111110111101111110111110001110111110111111111111111111001111111";
                    when "11001" => level_vec_out <= "1111110111101111110111111001110111110111111111111111111001111111";
                    when "11010" => level_vec_out <= "1111110111101111111111111001110111110111111111111111111001111111";
                    when "11011" => level_vec_out <= "1111110111101111111111111001110111110111111111111111111001111111";
                    when "11100" => level_vec_out <= "1111111111101111111111111101110111110111111111111111111001111111";
                    when "11101" => level_vec_out <= "1111111111111111111111111101111111110111111111111111111101111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111101111111110111111111111111111101111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111110111111111111111111101111111";
                when others => null;
                end case;
            when "101" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1011001100000001101101111111100010010101000101100110101111010111";
                    when "00001" => level_vec_out <= "1111001100000001101101111111111010010101000101100110101111010111";
                    when "00010" => level_vec_out <= "1111001100000001101101111111111010010101000101100110101111010111";
                    when "00011" => level_vec_out <= "1111001100000001101101111111111010010101001101100110101111010111";
                    when "00100" => level_vec_out <= "1111001110000001101101111111111010010101001101100110101111010111";
                    when "00101" => level_vec_out <= "1111001110010001101101111111111010010101001101100111101111010111";
                    when "00110" => level_vec_out <= "1111001110010001101101111111111010010101001101100111111111010111";
                    when "00111" => level_vec_out <= "1111001111110001101101111111111010010101001101100111111111010111";
                    when "01000" => level_vec_out <= "1111001111110001101101111111111010010101001101100111111111010111";
                    when "01001" => level_vec_out <= "1111001111110001111101111111111010010101001101100111111111010111";
                    when "01010" => level_vec_out <= "1111001111110001111101111111111010010101001101100111111111110111";
                    when "01011" => level_vec_out <= "1111101111110001111101111111111010010101001101100111111111110111";
                    when "01100" => level_vec_out <= "1111101111110001111101111111111010010101101101100111111111110111";
                    when "01101" => level_vec_out <= "1111101111110001111101111111111010010101101101100111111111110111";
                    when "01110" => level_vec_out <= "1111101111110001111101111111111110010101101101101111111111111111";
                    when "01111" => level_vec_out <= "1111101111110001111101111111111110010101101101101111111111111111";
                    when "10000" => level_vec_out <= "1111101111110001111101111111111110010101101101101111111111111111";
                    when "10001" => level_vec_out <= "1111101111110001111101111111111110010101101101101111111111111111";
                    when "10010" => level_vec_out <= "1111101111110001111101111111111110010101101101111111111111111111";
                    when "10011" => level_vec_out <= "1111101111110001111101111111111110010101101101111111111111111111";
                    when "10100" => level_vec_out <= "1111101111110101111101111111111110010111101101111111111111111111";
                    when "10101" => level_vec_out <= "1111101111110101111101111111111111010111101101111111111111111111";
                    when "10110" => level_vec_out <= "1111101111110101111101111111111111010111101101111111111111111111";
                    when "10111" => level_vec_out <= "1111101111110101111101111111111111010111101101111111111111111111";
                    when "11000" => level_vec_out <= "1111101111111101111101111111111111010111101101111111111111111111";
                    when "11001" => level_vec_out <= "1111101111111101111101111111111111111111101101111111111111111111";
                    when "11010" => level_vec_out <= "1111101111111101111101111111111111111111111111111111111111111111";
                    when "11011" => level_vec_out <= "1111101111111101111111111111111111111111111111111111111111111111";
                    when "11100" => level_vec_out <= "1111101111111111111111111111111111111111111111111111111111111111";
                    when "11101" => level_vec_out <= "1111101111111111111111111111111111111111111111111111111111111111";
                    when "11110" => level_vec_out <= "1111101111111111111111111111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111101111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "110" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0001111111111000111001111111011101110100110010101001100010001110";
                    when "00001" => level_vec_out <= "0001111111111000111001111111111101110101110010101001100010001110";
                    when "00010" => level_vec_out <= "0001111111111000111001111111111101110101110010101001100010001110";
                    when "00011" => level_vec_out <= "0001111111111000111001111111111101110101110010101001100010011111";
                    when "00100" => level_vec_out <= "0001111111111010111001111111111101110101110010101011100010011111";
                    when "00101" => level_vec_out <= "0001111111111010111001111111111101110101110011101011100010011111";
                    when "00110" => level_vec_out <= "0001111111111010111001111111111101110101110011101011100010011111";
                    when "00111" => level_vec_out <= "0001111111111010111001111111111101110101110011101011100010011111";
                    when "01000" => level_vec_out <= "0001111111111110111001111111111101110101110111101011100010011111";
                    when "01001" => level_vec_out <= "0001111111111110111101111111111101110101110111101011100010011111";
                    when "01010" => level_vec_out <= "0001111111111111111101111111111111110101110111101011100010011111";
                    when "01011" => level_vec_out <= "0001111111111111111101111111111111110111110111101011100010011111";
                    when "01100" => level_vec_out <= "0001111111111111111101111111111111110111110111101011100010011111";
                    when "01101" => level_vec_out <= "0101111111111111111101111111111111111111111111101011100010011111";
                    when "01110" => level_vec_out <= "0101111111111111111101111111111111111111111111101011100010011111";
                    when "01111" => level_vec_out <= "0101111111111111111101111111111111111111111111101011100110011111";
                    when "10000" => level_vec_out <= "0101111111111111111101111111111111111111111111101011100110011111";
                    when "10001" => level_vec_out <= "0101111111111111111101111111111111111111111111101011100110011111";
                    when "10010" => level_vec_out <= "0101111111111111111101111111111111111111111111101111100110011111";
                    when "10011" => level_vec_out <= "0101111111111111111101111111111111111111111111101111110110011111";
                    when "10100" => level_vec_out <= "0101111111111111111101111111111111111111111111101111110110011111";
                    when "10101" => level_vec_out <= "0101111111111111111101111111111111111111111111101111111110011111";
                    when "10110" => level_vec_out <= "0101111111111111111101111111111111111111111111101111111111111111";
                    when "10111" => level_vec_out <= "1111111111111111111101111111111111111111111111101111111111111111";
                    when "11000" => level_vec_out <= "1111111111111111111101111111111111111111111111101111111111111111";
                    when "11001" => level_vec_out <= "1111111111111111111101111111111111111111111111101111111111111111";
                    when "11010" => level_vec_out <= "1111111111111111111101111111111111111111111111101111111111111111";
                    when "11011" => level_vec_out <= "1111111111111111111101111111111111111111111111101111111111111111";
                    when "11100" => level_vec_out <= "1111111111111111111101111111111111111111111111101111111111111111";
                    when "11101" => level_vec_out <= "1111111111111111111101111111111111111111111111101111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111101111111111111111111111111101111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111101111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "111" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0000101101001010001100110110000000000110011000000011100111101010";
                    when "00001" => level_vec_out <= "0000101101001010001100110110000000000110011000000011100111101010";
                    when "00010" => level_vec_out <= "0000101101001010001100110110000010000110011000000111100111101010";
                    when "00011" => level_vec_out <= "0000101101001010001100110110000010000110011000000111100111101010";
                    when "00100" => level_vec_out <= "0000101101001010001100110110010010000110011000000111100111101010";
                    when "00101" => level_vec_out <= "0000111101001010001100110110010010000110111000000111100111101010";
                    when "00110" => level_vec_out <= "0000111101001010001100110110010010000110111000000111100111101010";
                    when "00111" => level_vec_out <= "0000111101011010001100110110010010000110111000000111100111101010";
                    when "01000" => level_vec_out <= "0000111101011010001100110110010010000110111000000111100111101010";
                    when "01001" => level_vec_out <= "0000111101011010001100110110010010000110111000000111100111101110";
                    when "01010" => level_vec_out <= "0000111101011010001100110110010010000111111000000111100111101110";
                    when "01011" => level_vec_out <= "0000111101011010001100110110010010010111111000000111100111101110";
                    when "01100" => level_vec_out <= "0000111101011010001100110110010010010111111000000111100111101110";
                    when "01101" => level_vec_out <= "1000111101011010001100110110011010010111111000000111101111101110";
                    when "01110" => level_vec_out <= "1000111101011010001100110110011010010111111000010111101111101110";
                    when "01111" => level_vec_out <= "1000111101011010001100110110011010010111111000010111101111101110";
                    when "10000" => level_vec_out <= "1000111101011010001100111110011010010111111000010111101111101110";
                    when "10001" => level_vec_out <= "1000111101011010001110111110111010010111111000010111101111101110";
                    when "10010" => level_vec_out <= "1000111101011010001110111110111010010111111000010111101111111110";
                    when "10011" => level_vec_out <= "1000111101011010001110111110111010110111111000010111101111111110";
                    when "10100" => level_vec_out <= "1000111101011010001110111110111010110111111001010111101111111110";
                    when "10101" => level_vec_out <= "1000111101011010001110111110111010110111111001010111101111111110";
                    when "10110" => level_vec_out <= "1000111101011010001110111110111010110111111001010111101111111110";
                    when "10111" => level_vec_out <= "1000111101011010101110111110111010110111111001010111101111111110";
                    when "11000" => level_vec_out <= "1010111111111010111110111110111010110111111001010111101111111110";
                    when "11001" => level_vec_out <= "1011111111111010111110111111111010110111111001010111101111111110";
                    when "11010" => level_vec_out <= "1111111111111010111110111111111010110111111001010111101111111110";
                    when "11011" => level_vec_out <= "1111111111111111111110111111111010110111111001010111101111111110";
                    when "11100" => level_vec_out <= "1111111111111111111110111111111010110111111001010111101111111111";
                    when "11101" => level_vec_out <= "1111111111111111111110111111111010110111111001011111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111011110111111101011111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when others => null;
        end case;
    end process;
end Behavioral;