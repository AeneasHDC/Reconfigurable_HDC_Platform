/**
 * @file level_hvec_gen_hdl.hpp
 * @brief This script generates HDL code for generating high-dimensional LEVEL vectors.
 * It is a novel method; for more information, please refer to our paper.
 *
 * @author Saeid Jamili and Marco Angioli
 * @note Author names are listed in alphabetical order.
 * @email <saeid.jamili@uniroma1.it>
 * @email <marco.angioli@uniroma1.it>
 *
 * @contributors
 *
 * @date Created: 24th July 2023
 * @date Last Updated: 23th August 2023
 *
 * @version 1.0.0
 *
 * @institute Sapienza University of Rome
 * @cite https://doi.org/10.xxxx/yyyyy
 *
 * @section DEPENDENCIES
 * - Dependency1: Description or version details.
 * - Dependency2: Description or version details.
 *
 * @section LICENSE
 * This file is part of the Aeneas HyperCompute Platform.
 *
 * Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 *
 * @section CHANGELOG
 * @version 1.0.0-dev - 23th August 2023
 * - Initial release
 *
 * @todo
 * - Complete level vector generator function
 * - Add training
 *
 * @see
 * -
 * -
 * -
 *
 */

module level_vec_gen (
    output reg [63:0] level_vec_out,
    input [2:0] frame_index,
    input [4:0] frame_id
);
    always @(*) begin
        // Update this function to match your requirements
        case (frame_index)
            0: begin
                case (frame_id)
                    0: level_vec_out = 64'b1100111111011010111110111111110001101110110100000001100111100101;
                    1: level_vec_out = 64'b1100111111011010111110111111110001101110110100000001100111100101;
                    2: level_vec_out = 64'b1100111111011010111110111111111001101110110110000001100111100101;
                    3: level_vec_out = 64'b1100111111011010111110111111111001101110110110010001100111100101;
                    4: level_vec_out = 64'b1100111111011010111110111111111101101110110110010001100111100101;
                    5: level_vec_out = 64'b1100111111011010111110111111111101101110110110011001100111100101;
                    6: level_vec_out = 64'b1100111111011010111110111111111101101110110110011001101111100101;
                    7: level_vec_out = 64'b1100111111011010111110111111111101101110110110011001101111100101;
                    8: level_vec_out = 64'b1100111111011010111110111111111101101110110110011001101111100101;
                    9: level_vec_out = 64'b1111111111011010111110111111111101101110110110011001101111100101;
                    10: level_vec_out = 64'b1111111111011010111110111111111101101110110110011001101111100101;
                    11: level_vec_out = 64'b1111111111011010111110111111111101101110110110011001101111100101;
                    12: level_vec_out = 64'b1111111111011010111110111111111101111110110110011001101111100101;
                    13: level_vec_out = 64'b1111111111011010111110111111111111111110110110011001101111100101;
                    14: level_vec_out = 64'b1111111111011010111110111111111111111110110110011001101111100101;
                    15: level_vec_out = 64'b1111111111011010111110111111111111111110110110011001101111100101;
                    16: level_vec_out = 64'b1111111111011010111110111111111111111110110110011011101111100101;
                    17: level_vec_out = 64'b1111111111011010111110111111111111111110111110011011101111100101;
                    18: level_vec_out = 64'b1111111111011010111110111111111111111110111110011011101111100111;
                    19: level_vec_out = 64'b1111111111011010111110111111111111111110111110011011101111100111;
                    20: level_vec_out = 64'b1111111111011010111110111111111111111110111110011011101111100111;
                    21: level_vec_out = 64'b1111111111011010111110111111111111111110111110011011101111100111;
                    22: level_vec_out = 64'b1111111111111010111110111111111111111110111111111111101111100111;
                    23: level_vec_out = 64'b1111111111111010111110111111111111111110111111111111101111100111;
                    24: level_vec_out = 64'b1111111111111010111110111111111111111110111111111111101111100111;
                    25: level_vec_out = 64'b1111111111111010111110111111111111111110111111111111101111101111;
                    26: level_vec_out = 64'b1111111111111110111111111111111111111111111111111111101111101111;
                    27: level_vec_out = 64'b1111111111111110111111111111111111111111111111111111101111101111;
                    28: level_vec_out = 64'b1111111111111110111111111111111111111111111111111111101111101111;
                    29: level_vec_out = 64'b1111111111111110111111111111111111111111111111111111101111101111;
                    30: level_vec_out = 64'b1111111111111110111111111111111111111111111111111111111111101111;
                    31: level_vec_out = 64'b1111111111111110111111111111111111111111111111111111111111101111;
                endcase
            end
            1: begin
                case (frame_id)
                    0: level_vec_out = 64'b1100011000111011100010011001100010000000100110010110000011010010;
                    1: level_vec_out = 64'b1100011000111011100010011001100010000000100110010110000011010010;
                    2: level_vec_out = 64'b1100011000111011100010011001100010000010100110010110000011010010;
                    3: level_vec_out = 64'b1100011000111011100010011001100010000010100110010110000011010010;
                    4: level_vec_out = 64'b1100011000111011100010011101100010000010100110010110100011010010;
                    5: level_vec_out = 64'b1100011000111011100010011101100010000010100110010111100011010010;
                    6: level_vec_out = 64'b1100011000111011100010011101100010000010100110010111100011010010;
                    7: level_vec_out = 64'b1100011000111011100010011101100010000011100110010111100011010010;
                    8: level_vec_out = 64'b1100011000111011100010011101100010000011100110010111100011110010;
                    9: level_vec_out = 64'b1100011000111011100010011101110010000011100110010111100011110010;
                    10: level_vec_out = 64'b1100011000111011100010011101110010000011100110010111100011110010;
                    11: level_vec_out = 64'b1100011000111011100010011101110010000011110110110111100011110110;
                    12: level_vec_out = 64'b1100011000111011100010011101110010000011110110110111100011110110;
                    13: level_vec_out = 64'b1110011000111011100010011101110010000011110110110111100011110110;
                    14: level_vec_out = 64'b1110011000111011100010011101110010000011110110110111100011110110;
                    15: level_vec_out = 64'b1110011000111011100010011101110010100011110110110111100011110111;
                    16: level_vec_out = 64'b1110011000111011100010011101110010100011110110110111100011110111;
                    17: level_vec_out = 64'b1110011100111011100010011101110010100011110110110111100011110111;
                    18: level_vec_out = 64'b1110011100111011100010011101110010100011110111110111100011110111;
                    19: level_vec_out = 64'b1110011100111011100010011101110011100011110111110111101011110111;
                    20: level_vec_out = 64'b1110011100111011100010011111110011100011110111111111101011110111;
                    21: level_vec_out = 64'b1110011101111011100010011111110011100011110111111111111011110111;
                    22: level_vec_out = 64'b1110011101111011100010011111110011100011110111111111111011110111;
                    23: level_vec_out = 64'b1110011101111011100010011111110011100011110111111111111011110111;
                    24: level_vec_out = 64'b1110011101111011100010011111110011100111111111111111111011110111;
                    25: level_vec_out = 64'b1110011101111011100010011111110111100111111111111111111011110111;
                    26: level_vec_out = 64'b1110011101111011100010011111110111101111111111111111111011110111;
                    27: level_vec_out = 64'b1110011101111011100011011111110111101111111111111111111011110111;
                    28: level_vec_out = 64'b1110011101111111101111111111110111101111111111111111111011111111;
                    29: level_vec_out = 64'b1111011101111111101111111111110111101111111111111111111011111111;
                    30: level_vec_out = 64'b1111111101111111111111111111111111101111111111111111111111111111;
                    31: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                endcase
            end
            2: begin
                case (frame_id)
                    0: level_vec_out = 64'b1101000011100001101001010111100001100100010001011011010011101110;
                    1: level_vec_out = 64'b1101000011100001101001010111100001100100010001011011010011101110;
                    2: level_vec_out = 64'b1101000011100001101001010111100001100100010001011011010011111110;
                    3: level_vec_out = 64'b1101000011100001111001010111100001100100010001011011010011111110;
                    4: level_vec_out = 64'b1101000011100001111001010111100001100100010011011011010011111110;
                    5: level_vec_out = 64'b1101000011100001111001010111100001100100010011011011010011111110;
                    6: level_vec_out = 64'b1101000011100001111001010111100001100100010011011011010011111110;
                    7: level_vec_out = 64'b1101000011100001111001010111100001100100010011011011010011111110;
                    8: level_vec_out = 64'b1101000011100001111001010111100001100110010011011011010011111110;
                    9: level_vec_out = 64'b1101010011100001111001010111100001100110010011011011010011111110;
                    10: level_vec_out = 64'b1101010011100001111001010111100001110111010011011011010011111110;
                    11: level_vec_out = 64'b1101010011100001111001110111100001110111010011011011010011111110;
                    12: level_vec_out = 64'b1101011011100101111001110111100001110111010011111011010011111110;
                    13: level_vec_out = 64'b1101011011100101111001110111100011110111010011111011010011111110;
                    14: level_vec_out = 64'b1101011011100101111001110111100011110111010011111011010011111111;
                    15: level_vec_out = 64'b1101011011100101111001110111100011110111010011111111010011111111;
                    16: level_vec_out = 64'b1101011011100101111001110111100011111111010011111111010011111111;
                    17: level_vec_out = 64'b1101011111100101111001110111101011111111010011111111010011111111;
                    18: level_vec_out = 64'b1101011111100101111101110111101011111111010011111111010011111111;
                    19: level_vec_out = 64'b1101011111100101111111111111101011111111010011111111010011111111;
                    20: level_vec_out = 64'b1101011111100101111111111111101011111111010011111111010011111111;
                    21: level_vec_out = 64'b1101011111100101111111111111101011111111011011111111010011111111;
                    22: level_vec_out = 64'b1101011111100101111111111111101011111111011011111111010011111111;
                    23: level_vec_out = 64'b1101011111100101111111111111111011111111011011111111010011111111;
                    24: level_vec_out = 64'b1101111111100101111111111111111011111111011011111111011011111111;
                    25: level_vec_out = 64'b1101111111100101111111111111111111111111011011111111011011111111;
                    26: level_vec_out = 64'b1101111111100101111111111111111111111111011011111111111011111111;
                    27: level_vec_out = 64'b1101111111110101111111111111111111111111111011111111111011111111;
                    28: level_vec_out = 64'b1101111111110101111111111111111111111111111011111111111011111111;
                    29: level_vec_out = 64'b1101111111110101111111111111111111111111111111111111111011111111;
                    30: level_vec_out = 64'b1101111111110101111111111111111111111111111111111111111011111111;
                    31: level_vec_out = 64'b1111111111111101111111111111111111111111111111111111111111111111;
                endcase
            end
            3: begin
                case (frame_id)
                    0: level_vec_out = 64'b0111110001001110101001000111100111000101101010000101100111110101;
                    1: level_vec_out = 64'b0111110101001110101001000111101111000101101010000101100111111101;
                    2: level_vec_out = 64'b0111110101001110101001000111101111000101101010000101100111111101;
                    3: level_vec_out = 64'b0111110101001110101001000111101111000101101010000101100111111101;
                    4: level_vec_out = 64'b0111110101001110101001000111101111000111111010000101100111111101;
                    5: level_vec_out = 64'b0111110101001110101001000111101111000111111010000101100111111101;
                    6: level_vec_out = 64'b0111110101001110101001000111101111000111111010000101100111111111;
                    7: level_vec_out = 64'b0111110101001110101011000111101111000111111010000111100111111111;
                    8: level_vec_out = 64'b0111110101001110101011000111101111000111111010000111100111111111;
                    9: level_vec_out = 64'b0111110101001110101011010111101111000111111010000111100111111111;
                    10: level_vec_out = 64'b0111110101001110101011010111101111000111111010000111101111111111;
                    11: level_vec_out = 64'b0111110101001110101011010111101111000111111010000111101111111111;
                    12: level_vec_out = 64'b0111110101001110101011010111101111000111111010000111101111111111;
                    13: level_vec_out = 64'b0111110101001110101011010111111111000111111010000111101111111111;
                    14: level_vec_out = 64'b0111110101001110101011010111111111100111111110000111101111111111;
                    15: level_vec_out = 64'b0111110101001110101011010111111111100111111110100111101111111111;
                    16: level_vec_out = 64'b0111110101001110101011010111111111100111111110100111101111111111;
                    17: level_vec_out = 64'b0111110111001110101011011111111111100111111110100111101111111111;
                    18: level_vec_out = 64'b0111110111001110111011011111111111100111111110110111101111111111;
                    19: level_vec_out = 64'b0111110111001110111011011111111111100111111110110111101111111111;
                    20: level_vec_out = 64'b0111110111011110111011011111111111100111111110110111101111111111;
                    21: level_vec_out = 64'b0111110111011110111011011111111111100111111110110111101111111111;
                    22: level_vec_out = 64'b1111110111011110111011011111111111100111111110110111101111111111;
                    23: level_vec_out = 64'b1111110111011110111111011111111111100111111110110111101111111111;
                    24: level_vec_out = 64'b1111110111011110111111011111111111110111111110110111101111111111;
                    25: level_vec_out = 64'b1111110111011111111111011111111111110111111110110111101111111111;
                    26: level_vec_out = 64'b1111110111011111111111011111111111110111111110110111101111111111;
                    27: level_vec_out = 64'b1111110111011111111111111111111111110111111110111111101111111111;
                    28: level_vec_out = 64'b1111110111011111111111111111111111110111111110111111101111111111;
                    29: level_vec_out = 64'b1111110111011111111111111111111111111111111110111111111111111111;
                    30: level_vec_out = 64'b1111110111011111111111111111111111111111111111111111111111111111;
                    31: level_vec_out = 64'b1111111111011111111111111111111111111111111111111111111111111111;
                endcase
            end
            4: begin
                case (frame_id)
                    0: level_vec_out = 64'b1011101111001001001011101110001101100100001100110001110010101011;
                    1: level_vec_out = 64'b1011101111001001001011101110001101100100001100110001110010101011;
                    2: level_vec_out = 64'b1011101111001001101011101110001101100100001100110001110010101011;
                    3: level_vec_out = 64'b1011101111001001101011101110001101100100001100110001110010101011;
                    4: level_vec_out = 64'b1011101111001001101111101110001101100100001100110001110010111011;
                    5: level_vec_out = 64'b1011101111001001101111101110001101100100001100110101110010111011;
                    6: level_vec_out = 64'b1011101111001001101111101110001101100110001100110101110010111011;
                    7: level_vec_out = 64'b1011101111001001101111101110001101100110001100110101110010111011;
                    8: level_vec_out = 64'b1011101111001011101111101110001111100110011100110101110010111011;
                    9: level_vec_out = 64'b1011101111001011101111101110001111100110011110110111110010111011;
                    10: level_vec_out = 64'b1011101111001011101111101110101111100110011110110111110011111111;
                    11: level_vec_out = 64'b1011101111001011101111101110101111100110011110110111111011111111;
                    12: level_vec_out = 64'b1011101111001011101111101110101111100110011110110111111011111111;
                    13: level_vec_out = 64'b1011101111001011111111101110101111110111011110110111111011111111;
                    14: level_vec_out = 64'b1011101111001011111111101110101111111111011110110111111011111111;
                    15: level_vec_out = 64'b1011101111001011111111101110101111111111011110111111111011111111;
                    16: level_vec_out = 64'b1011111111101011111111101110101111111111011110111111111011111111;
                    17: level_vec_out = 64'b1011111111101011111111101110101111111111011110111111111011111111;
                    18: level_vec_out = 64'b1011111111101011111111101110101111111111011110111111111011111111;
                    19: level_vec_out = 64'b1011111111101011111111101110101111111111011110111111111011111111;
                    20: level_vec_out = 64'b1011111111101111111111101110101111111111011110111111111011111111;
                    21: level_vec_out = 64'b1011111111101111111111101110101111111111011110111111111011111111;
                    22: level_vec_out = 64'b1111111111101111111111101110101111111111011110111111111011111111;
                    23: level_vec_out = 64'b1111111111101111111111101110101111111111111110111111111011111111;
                    24: level_vec_out = 64'b1111111111101111111111101111101111111111111110111111111011111111;
                    25: level_vec_out = 64'b1111111111101111111111101111101111111111111110111111111011111111;
                    26: level_vec_out = 64'b1111111111101111111111101111101111111111111110111111111111111111;
                    27: level_vec_out = 64'b1111111111101111111111101111111111111111111110111111111111111111;
                    28: level_vec_out = 64'b1111111111101111111111101111111111111111111110111111111111111111;
                    29: level_vec_out = 64'b1111111111101111111111111111111111111111111111111111111111111111;
                    30: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    31: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                endcase
            end
            5: begin
                case (frame_id)
                    0: level_vec_out = 64'b1110100110001001101011100011110010101110001000110100001100110010;
                    1: level_vec_out = 64'b1110100110001001101111110011110010111110001100110100001100110010;
                    2: level_vec_out = 64'b1110100110001001101111110011110010111110001100110100001100110010;
                    3: level_vec_out = 64'b1110100110001101101111110011110010111110001100110100001100110010;
                    4: level_vec_out = 64'b1110100110001101101111110011110010111110001100110100001100110010;
                    5: level_vec_out = 64'b1110100110001101101111110011111010111110001100110100001100110010;
                    6: level_vec_out = 64'b1110100110001101101111110011111110111110001100110100001100110010;
                    7: level_vec_out = 64'b1111100110001101101111110011111110111110001100110110001110110110;
                    8: level_vec_out = 64'b1111100110001101101111110011111110111110001100110110001110110110;
                    9: level_vec_out = 64'b1111100110001101101111110011111110111110001100110110001110110110;
                    10: level_vec_out = 64'b1111100110001101101111110011111110111110001100110110001110110110;
                    11: level_vec_out = 64'b1111100110001101101111111011111110111110001100110110001110110110;
                    12: level_vec_out = 64'b1111100111001101101111111011111110111110001100110110001110110110;
                    13: level_vec_out = 64'b1111100111001101101111111011111110111110001100110110001110110110;
                    14: level_vec_out = 64'b1111100111001101101111111011111110111110011100110110001111110110;
                    15: level_vec_out = 64'b1111100111001101101111111011111110111110011100110110001111110110;
                    16: level_vec_out = 64'b1111100111001111101111111011111110111110011100110110001111110110;
                    17: level_vec_out = 64'b1111100111001111101111111011111111111110011100110110001111111110;
                    18: level_vec_out = 64'b1111100111001111101111111011111111111110011100110110101111111110;
                    19: level_vec_out = 64'b1111101111101111101111111011111111111110011100110110101111111110;
                    20: level_vec_out = 64'b1111101111101111101111111011111111111110011100110110101111111110;
                    21: level_vec_out = 64'b1111101111111111101111111011111111111110011101110111101111111110;
                    22: level_vec_out = 64'b1111101111111111111111111011111111111110011101110111101111111110;
                    23: level_vec_out = 64'b1111101111111111111111111011111111111110111101110111101111111110;
                    24: level_vec_out = 64'b1111101111111111111111111011111111111110111101110111101111111110;
                    25: level_vec_out = 64'b1111111111111111111111111011111111111110111111110111101111111110;
                    26: level_vec_out = 64'b1111111111111111111111111011111111111110111111111111101111111110;
                    27: level_vec_out = 64'b1111111111111111111111111011111111111111111111111111101111111110;
                    28: level_vec_out = 64'b1111111111111111111111111011111111111111111111111111101111111111;
                    29: level_vec_out = 64'b1111111111111111111111111011111111111111111111111111101111111111;
                    30: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111101111111111;
                    31: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                endcase
            end
            6: begin
                case (frame_id)
                    0: level_vec_out = 64'b0010100000111000100101111101010010011010011100100010100111110010;
                    1: level_vec_out = 64'b0010100001111000100101111101010010011010011100100010100111110010;
                    2: level_vec_out = 64'b0010101001111000100101111101010010011010011100100010100111110010;
                    3: level_vec_out = 64'b0010111001111000110101111101010010011010011100100011100111110011;
                    4: level_vec_out = 64'b0010111001111000110101111101010010011010011100100011100111110011;
                    5: level_vec_out = 64'b0010111001111100110101111111010010011010011100100011100111110011;
                    6: level_vec_out = 64'b1010111001111100110101111111010010011010011110100011110111110011;
                    7: level_vec_out = 64'b1010111001111100110101111111010010011110011110100011110111110011;
                    8: level_vec_out = 64'b1010111001111100110101111111010010011110011110100011110111110011;
                    9: level_vec_out = 64'b1010111001111100110101111111010010011110011110100011110111110011;
                    10: level_vec_out = 64'b1010111001111100110101111111010010011110011110100011110111110011;
                    11: level_vec_out = 64'b1010111001111100110101111111010010011110011110100011110111110011;
                    12: level_vec_out = 64'b1011111001111101110101111111010010111110011110100011110111110011;
                    13: level_vec_out = 64'b1011111001111111110101111111010010111110011110100011110111110011;
                    14: level_vec_out = 64'b1011111001111111110101111111011010111110111110100011110111110011;
                    15: level_vec_out = 64'b1011111001111111110101111111011010111110111110100011110111110011;
                    16: level_vec_out = 64'b1111111011111111110101111111011010111110111110100011110111110011;
                    17: level_vec_out = 64'b1111111011111111110101111111011010111110111110100011110111110011;
                    18: level_vec_out = 64'b1111111011111111110101111111011010111110111110101011110111110011;
                    19: level_vec_out = 64'b1111111011111111110101111111011010111110111110101011110111110011;
                    20: level_vec_out = 64'b1111111111111111110101111111011010111110111111101011110111110011;
                    21: level_vec_out = 64'b1111111111111111110101111111011010111110111111101011110111111011;
                    22: level_vec_out = 64'b1111111111111111110101111111011010111110111111101011111111111011;
                    23: level_vec_out = 64'b1111111111111111110101111111111011111111111111101011111111111111;
                    24: level_vec_out = 64'b1111111111111111110101111111111011111111111111101011111111111111;
                    25: level_vec_out = 64'b1111111111111111110101111111111011111111111111101011111111111111;
                    26: level_vec_out = 64'b1111111111111111110101111111111011111111111111101011111111111111;
                    27: level_vec_out = 64'b1111111111111111110111111111111011111111111111101011111111111111;
                    28: level_vec_out = 64'b1111111111111111111111111111111011111111111111101011111111111111;
                    29: level_vec_out = 64'b1111111111111111111111111111111011111111111111111011111111111111;
                    30: level_vec_out = 64'b1111111111111111111111111111111011111111111111111011111111111111;
                    31: level_vec_out = 64'b1111111111111111111111111111111011111111111111111011111111111111;
                endcase
            end
            7: begin
                case (frame_id)
                    0: level_vec_out = 64'b1010000011110010010001101000011111100111001000100101011000101110;
                    1: level_vec_out = 64'b1010000011110010010001101000011111100111001000100101011000101110;
                    2: level_vec_out = 64'b1010100011110010010001101000011111100111001000101101011000101110;
                    3: level_vec_out = 64'b1010100011110010010001101000011111100111001000101101011000111110;
                    4: level_vec_out = 64'b1010100011110010010001101000011111100111001000101101011000111110;
                    5: level_vec_out = 64'b1010100011110010010001101100011111100111001000101111011000111110;
                    6: level_vec_out = 64'b1010100111110010010001101100011111100111001000101111011000111110;
                    7: level_vec_out = 64'b1010100111110010010001101100011111100111001000101111011000111110;
                    8: level_vec_out = 64'b1011100111110010010001101100011111100111001100101111111000111110;
                    9: level_vec_out = 64'b1011100111110010010001101101011111100111001100101111111000111110;
                    10: level_vec_out = 64'b1011100111110010010001101101111111100111001100101111111010111110;
                    11: level_vec_out = 64'b1011100111110010010101101101111111100111001100101111111011111110;
                    12: level_vec_out = 64'b1011100111110010010101101101111111100111001100101111111011111110;
                    13: level_vec_out = 64'b1011100111110010010101101101111111100111001100101111111011111110;
                    14: level_vec_out = 64'b1011100111110010010101101101111111100111001100101111111011111110;
                    15: level_vec_out = 64'b1011100111110010011101101111111111110111001100101111111011111110;
                    16: level_vec_out = 64'b1011100111110010011101101111111111111111001100101111111011111110;
                    17: level_vec_out = 64'b1011100111110010011101101111111111111111001100101111111011111110;
                    18: level_vec_out = 64'b1011100111110010011111101111111111111111001100101111111011111110;
                    19: level_vec_out = 64'b1011100111110011011111101111111111111111001101101111111011111110;
                    20: level_vec_out = 64'b1011110111110011011111101111111111111111101101101111111011111110;
                    21: level_vec_out = 64'b1011110111110011111111101111111111111111101101101111111011111110;
                    22: level_vec_out = 64'b1011110111110011111111101111111111111111101101101111111011111110;
                    23: level_vec_out = 64'b1011110111110011111111101111111111111111101101101111111011111110;
                    24: level_vec_out = 64'b1111110111110011111111111111111111111111101101101111111011111110;
                    25: level_vec_out = 64'b1111110111110011111111111111111111111111101111111111111011111110;
                    26: level_vec_out = 64'b1111110111110011111111111111111111111111101111111111111111111110;
                    27: level_vec_out = 64'b1111110111110011111111111111111111111111101111111111111111111110;
                    28: level_vec_out = 64'b1111110111110011111111111111111111111111111111111111111111111110;
                    29: level_vec_out = 64'b1111110111110111111111111111111111111111111111111111111111111110;
                    30: level_vec_out = 64'b1111110111110111111111111111111111111111111111111111111111111110;
                    31: level_vec_out = 64'b1111110111110111111111111111111111111111111111111111111111111111;
                endcase
            end
        endcase
    end
endmodule