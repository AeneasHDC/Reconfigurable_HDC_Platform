/**
 * @file level_hvec_gen_hdl.hpp
 * @brief This script generates HDL code for generating high-dimensional LEVEL vectors.
 * It is a novel method; for more information, please refer to our paper.
 *
 * @author Saeid Jamili and Marco Angioli
 * @note Author names are listed in alphabetical order.
 * @email <saeid.jamili@uniroma1.it>
 * @email <marco.angioli@uniroma1.it>
 *
 * @contributors
 *
 * @date Created: 24th July 2023
 * @date Last Updated: 23th August 2023
 *
 * @version 1.0.0
 *
 * @institute Sapienza University of Rome
 * @cite https://doi.org/10.xxxx/yyyyy
 *
 * @section DEPENDENCIES
 * - Dependency1: Description or version details.
 * - Dependency2: Description or version details.
 *
 * @section LICENSE
 * This file is part of the Aeneas HyperCompute Platform.
 *
 * Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 *
 * @section CHANGELOG
 * @version 1.0.0-dev - 23th August 2023
 * - Initial release
 *
 * @todo
 * - Complete level vector generator function
 * - Add training
 *
 * @see
 * -
 * -
 * -
 *
 */

module level_hvec_gen #(parameter int DI_PARALLEL_W_BITS = 64) (
  input logic [2:0] frame_index,
  input logic [4:0] frame_id,
  output logic [DI_PARALLEL_W_BITS-1:0] level_vec_out
);
  always_comb begin
    case (frame_index)
      0:
        case (frame_id)
          0:
            level_vec_out = 64'b1110010100010001000010111001100101010000011000000101100100101110;
          1:
            level_vec_out = 64'b1110010110010001000010111001100101011000011000000101100100101110;
          2:
            level_vec_out = 64'b1110010111010011000010111001100101011000011000000101100100101110;
          3:
            level_vec_out = 64'b1110010111010011000010111001100101011000011000000101100100101110;
          4:
            level_vec_out = 64'b1110010111010011000010111001100101011000011000100101100100101110;
          5:
            level_vec_out = 64'b1110010111010011000010111001100101011000011000100101100100101110;
          6:
            level_vec_out = 64'b1110010111010011000010111001101101011000011000100101100100111110;
          7:
            level_vec_out = 64'b1110010111011011000010111001101111011000011000100101100100111110;
          8:
            level_vec_out = 64'b1110010111011011000010111001101111011000011000100101100100111110;
          9:
            level_vec_out = 64'b1110010111011011000010111001111111011000011000100101100100111110;
          10:
            level_vec_out = 64'b1110010111011011000010111001111111011000011000100101100100111110;
          11:
            level_vec_out = 64'b1110010111011011000010111001111111011000011000100101100100111110;
          12:
            level_vec_out = 64'b1110010111011011100010111001111111011001011010100101100100111110;
          13:
            level_vec_out = 64'b1110011111011011100010111011111111011001011010100101100100111110;
          14:
            level_vec_out = 64'b1111011111011011100010111011111111011001111111100111100100111110;
          15:
            level_vec_out = 64'b1111011111011011101010111011111111111001111111100111100100111110;
          16:
            level_vec_out = 64'b1111011111011011101010111011111111111001111111100111100100111110;
          17:
            level_vec_out = 64'b1111011111011011111010111011111111111001111111100111100101111110;
          18:
            level_vec_out = 64'b1111011111011111111010111011111111111001111111101111100111111110;
          19:
            level_vec_out = 64'b1111011111011111111110111011111111111001111111101111100111111110;
          20:
            level_vec_out = 64'b1111011111011111111110111111111111111011111111101111110111111110;
          21:
            level_vec_out = 64'b1111011111011111111111111111111111111011111111101111110111111110;
          22:
            level_vec_out = 64'b1111011111011111111111111111111111111011111111101111110111111110;
          23:
            level_vec_out = 64'b1111011111011111111111111111111111111011111111101111110111111110;
          24:
            level_vec_out = 64'b1111011111011111111111111111111111111011111111101111110111111110;
          25:
            level_vec_out = 64'b1111011111011111111111111111111111111011111111101111110111111110;
          26:
            level_vec_out = 64'b1111011111011111111111111111111111111011111111101111110111111110;
          27:
            level_vec_out = 64'b1111011111011111111111111111111111111011111111101111110111111110;
          28:
            level_vec_out = 64'b1111011111011111111111111111111111111011111111101111110111111111;
          29:
            level_vec_out = 64'b1111011111011111111111111111111111111111111111101111110111111111;
          30:
            level_vec_out = 64'b1111111111011111111111111111111111111111111111101111111111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111101111111111111111;
        endcase
      1:
        case (frame_id)
          0:
            level_vec_out = 64'b0010110111110111011111001100111101111010110011101101000110000100;
          1:
            level_vec_out = 64'b1010110111110111011111001100111101111010110011101101000110000100;
          2:
            level_vec_out = 64'b1010110111110111011111001100111101111010110011101101000110000100;
          3:
            level_vec_out = 64'b1010110111110111011111001100111101111010110011101101000110000100;
          4:
            level_vec_out = 64'b1010110111110111011111001100111101111010110011101101000110000100;
          5:
            level_vec_out = 64'b1010110111110111011111001100111101111010110011111101000110000100;
          6:
            level_vec_out = 64'b1010110111110111011111001100111111111010110011111101000110000100;
          7:
            level_vec_out = 64'b1010110111110111011111001100111111111010110011111101000110000100;
          8:
            level_vec_out = 64'b1010110111110111011111001100111111111010110111111101100110001100;
          9:
            level_vec_out = 64'b1010110111110111011111001100111111111010110111111101100110001100;
          10:
            level_vec_out = 64'b1010110111110111011111001110111111111010110111111101100110001100;
          11:
            level_vec_out = 64'b1010110111110111011111001110111111111110110111111101100110001100;
          12:
            level_vec_out = 64'b1010110111110111011111001110111111111110110111111101100110001100;
          13:
            level_vec_out = 64'b1010110111110111011111001110111111111110110111111101100110001100;
          14:
            level_vec_out = 64'b1010110111110111011111001110111111111110110111111101100110001100;
          15:
            level_vec_out = 64'b1010110111110111011111011110111111111110110111111101100110001100;
          16:
            level_vec_out = 64'b1010110111110111011111011110111111111110110111111101100110001100;
          17:
            level_vec_out = 64'b1110110111110111011111111110111111111110110111111101100110001110;
          18:
            level_vec_out = 64'b1110110111110111011111111110111111111110110111111101100110001110;
          19:
            level_vec_out = 64'b1110110111110111011111111110111111111110110111111101100110011110;
          20:
            level_vec_out = 64'b1110110111110111011111111110111111111110110111111101100110011110;
          21:
            level_vec_out = 64'b1110110111110111011111111110111111111111110111111101100110011110;
          22:
            level_vec_out = 64'b1110110111110111011111111110111111111111110111111101100110011111;
          23:
            level_vec_out = 64'b1110110111111111011111111110111111111111110111111101100110011111;
          24:
            level_vec_out = 64'b1110110111111111111111111110111111111111111111111101100110011111;
          25:
            level_vec_out = 64'b1111110111111111111111111110111111111111111111111101110110011111;
          26:
            level_vec_out = 64'b1111110111111111111111111110111111111111111111111101110110111111;
          27:
            level_vec_out = 64'b1111110111111111111111111110111111111111111111111101110111111111;
          28:
            level_vec_out = 64'b1111110111111111111111111110111111111111111111111101110111111111;
          29:
            level_vec_out = 64'b1111110111111111111111111110111111111111111111111101110111111111;
          30:
            level_vec_out = 64'b1111111111111111111111111110111111111111111111111101110111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111101110111111111;
        endcase
      2:
        case (frame_id)
          0:
            level_vec_out = 64'b1000111101110111010000010011000001010110110000101101000001100010;
          1:
            level_vec_out = 64'b1000111101110111010000010011000001010110110000101101001001100010;
          2:
            level_vec_out = 64'b1000111101110111010000010011100001010110110000101101001001100010;
          3:
            level_vec_out = 64'b1000111101110111010000010011100001110110110000101101101001100010;
          4:
            level_vec_out = 64'b1000111101110111010000010011100001110110110000101101101001100010;
          5:
            level_vec_out = 64'b1000111101110111010000010011100001110110110001101101101001100010;
          6:
            level_vec_out = 64'b1000111101110111110010010011100011110110110001101101101001100010;
          7:
            level_vec_out = 64'b1000111101110111110010010011100011110110110001101101101001100010;
          8:
            level_vec_out = 64'b1000111101110111110010010011101011110110110011101101101001100010;
          9:
            level_vec_out = 64'b1000111101110111110010010011101011110110110011101101101001100010;
          10:
            level_vec_out = 64'b1000111101110111110010010011101011110110110011101101101001100010;
          11:
            level_vec_out = 64'b1000111101110111110010010011101011110110110011101101101001100010;
          12:
            level_vec_out = 64'b1000111101110111110010010111101011111110110011101101101001100010;
          13:
            level_vec_out = 64'b1000111101110111111010010111101011111110110011101101101001100010;
          14:
            level_vec_out = 64'b1000111101110111111010010111101011111110110111101101101001100010;
          15:
            level_vec_out = 64'b1000111101110111111010010111101011111110110111101101101011100010;
          16:
            level_vec_out = 64'b1000111101110111111010010111101011111110110111101101101011100010;
          17:
            level_vec_out = 64'b1000111101110111111010010111101011111110110111101101101011100010;
          18:
            level_vec_out = 64'b1000111111110111111010010111101011111110110111101101101011100010;
          19:
            level_vec_out = 64'b1000111111110111111010010111101111111110110111101101101111100010;
          20:
            level_vec_out = 64'b1001111111110111111110110111101111111110110111101101101111100010;
          21:
            level_vec_out = 64'b1001111111110111111110111111101111111110110111101101101111100011;
          22:
            level_vec_out = 64'b1001111111111111111110111111101111111110110111111101101111100011;
          23:
            level_vec_out = 64'b1001111111111111111110111111101111111110110111111101101111100011;
          24:
            level_vec_out = 64'b1001111111111111111110111111101111111110110111111101101111100011;
          25:
            level_vec_out = 64'b1001111111111111111110111111101111111110110111111101101111101111;
          26:
            level_vec_out = 64'b1101111111111111111111111111101111111110110111111101101111101111;
          27:
            level_vec_out = 64'b1101111111111111111111111111101111111111110111111101101111101111;
          28:
            level_vec_out = 64'b1101111111111111111111111111101111111111111111111101111111111111;
          29:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111101111111111111;
          30:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        endcase
      3:
        case (frame_id)
          0:
            level_vec_out = 64'b1101000111010111010100100011110011010010001001100001000111111110;
          1:
            level_vec_out = 64'b1101000111010111010100110011110011010010001001100001000111111110;
          2:
            level_vec_out = 64'b1101000111010111010100110011110011010010001001100001000111111110;
          3:
            level_vec_out = 64'b1101000111010111010100110011110011010010001001100011000111111110;
          4:
            level_vec_out = 64'b1101000111010111010100110011110011010010001001100011000111111110;
          5:
            level_vec_out = 64'b1101101111010111010110110011110011010010001011100011000111111110;
          6:
            level_vec_out = 64'b1101101111010111010110110011110011010010001011100011000111111110;
          7:
            level_vec_out = 64'b1101101111010111010110110111110011010010001011100011000111111110;
          8:
            level_vec_out = 64'b1101101111010111010110110111110011010010001011100011000111111110;
          9:
            level_vec_out = 64'b1101101111010111010110111111110011010010001011100011000111111111;
          10:
            level_vec_out = 64'b1101111111010111010110111111110011010010001011100011000111111111;
          11:
            level_vec_out = 64'b1101111111010111010110111111110011010010001011100011000111111111;
          12:
            level_vec_out = 64'b1101111111010111010110111111110011010010001011100011000111111111;
          13:
            level_vec_out = 64'b1101111111010111010110111111110011010010011011100011100111111111;
          14:
            level_vec_out = 64'b1101111111010111010110111111110011010010011011100011100111111111;
          15:
            level_vec_out = 64'b1101111111010111010110111111110011010010111011100111100111111111;
          16:
            level_vec_out = 64'b1101111111010111010110111111110011010011111011100111101111111111;
          17:
            level_vec_out = 64'b1101111111010111010111111111110011010011111011100111101111111111;
          18:
            level_vec_out = 64'b1101111111010111010111111111110011011011111011100111101111111111;
          19:
            level_vec_out = 64'b1101111111010111010111111111110011011011111111100111101111111111;
          20:
            level_vec_out = 64'b1101111111010111010111111111110011011011111111100111101111111111;
          21:
            level_vec_out = 64'b1101111111010111010111111111110011011011111111100111101111111111;
          22:
            level_vec_out = 64'b1101111111111111110111111111110011011011111111100111101111111111;
          23:
            level_vec_out = 64'b1101111111111111110111111111110011011011111111100111101111111111;
          24:
            level_vec_out = 64'b1101111111111111110111111111110011011011111111100111101111111111;
          25:
            level_vec_out = 64'b1101111111111111110111111111110011011011111111100111101111111111;
          26:
            level_vec_out = 64'b1101111111111111110111111111110011011111111111100111101111111111;
          27:
            level_vec_out = 64'b1101111111111111110111111111110011011111111111110111101111111111;
          28:
            level_vec_out = 64'b1101111111111111110111111111110011111111111111110111101111111111;
          29:
            level_vec_out = 64'b1111111111111111111111111111110011111111111111110111111111111111;
          30:
            level_vec_out = 64'b1111111111111111111111111111110111111111111111110111111111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111110111111111111111111111111111111111;
        endcase
      4:
        case (frame_id)
          0:
            level_vec_out = 64'b1001010010101000101101001011011101110001111111100011000001001111;
          1:
            level_vec_out = 64'b1001010010101000101101001011011101110001111111100011000001001111;
          2:
            level_vec_out = 64'b1001010110101000101101001011011101110001111111100011000001001111;
          3:
            level_vec_out = 64'b1001010110101000101101001011011101110001111111100011000001001111;
          4:
            level_vec_out = 64'b1001010110101000101101001011011101110001111111100011000001001111;
          5:
            level_vec_out = 64'b1001010110101000101101001011011101110001111111100011000001011111;
          6:
            level_vec_out = 64'b1001010110101000101111001011011101110001111111100011000001011111;
          7:
            level_vec_out = 64'b1001010110101000101111001011011101111001111111100011000001011111;
          8:
            level_vec_out = 64'b1001010110101000101111001011011101111001111111100011000001111111;
          9:
            level_vec_out = 64'b1001010110101000101111001011011101111001111111101011000001111111;
          10:
            level_vec_out = 64'b1001011110101001101111001011011101111001111111101011000001111111;
          11:
            level_vec_out = 64'b1001011110101001101111001011011101111001111111101011000001111111;
          12:
            level_vec_out = 64'b1001011110101001101111001011011101111001111111101011000001111111;
          13:
            level_vec_out = 64'b1001011110101001101111001011011101111001111111101111000001111111;
          14:
            level_vec_out = 64'b1101011110101001101111001111011101111001111111101111000001111111;
          15:
            level_vec_out = 64'b1111011110101001111111001111011101111001111111101111000001111111;
          16:
            level_vec_out = 64'b1111011110101111111111001111011101111001111111101111000001111111;
          17:
            level_vec_out = 64'b1111011110101111111111001111011101111001111111101111000001111111;
          18:
            level_vec_out = 64'b1111011110101111111111001111011101111001111111101111000001111111;
          19:
            level_vec_out = 64'b1111111110101111111111001111011101111011111111101111000011111111;
          20:
            level_vec_out = 64'b1111111110101111111111001111011101111011111111101111000011111111;
          21:
            level_vec_out = 64'b1111111110101111111111101111011101111011111111101111000011111111;
          22:
            level_vec_out = 64'b1111111110101111111111101111011101111011111111101111000011111111;
          23:
            level_vec_out = 64'b1111111110101111111111101111011101111011111111111111000011111111;
          24:
            level_vec_out = 64'b1111111110101111111111101111011101111111111111111111000111111111;
          25:
            level_vec_out = 64'b1111111110101111111111101111011101111111111111111111000111111111;
          26:
            level_vec_out = 64'b1111111110101111111111101111111101111111111111111111100111111111;
          27:
            level_vec_out = 64'b1111111110101111111111101111111101111111111111111111101111111111;
          28:
            level_vec_out = 64'b1111111110101111111111101111111101111111111111111111101111111111;
          29:
            level_vec_out = 64'b1111111110101111111111101111111101111111111111111111101111111111;
          30:
            level_vec_out = 64'b1111111111101111111111101111111101111111111111111111101111111111;
          31:
            level_vec_out = 64'b1111111111101111111111101111111101111111111111111111111111111111;
        endcase
      5:
        case (frame_id)
          0:
            level_vec_out = 64'b0011011101011000000001110100100101111110111011110101001100101011;
          1:
            level_vec_out = 64'b0011011101011000000001110100100101111110111011110101001110101011;
          2:
            level_vec_out = 64'b0011011101011001000001110101100101111110111011110101001110101011;
          3:
            level_vec_out = 64'b0111011101011101000001110111100101111110111011110101001110101011;
          4:
            level_vec_out = 64'b0111011101011101000001110111100101111110111011110101001110101011;
          5:
            level_vec_out = 64'b0111011101011111000001110111100101111110111011110101001110101011;
          6:
            level_vec_out = 64'b0111011101011111000001110111100101111110111011110101001110101011;
          7:
            level_vec_out = 64'b0111011101011111000001110111101101111110111011110101001110101011;
          8:
            level_vec_out = 64'b0111011111011111000001110111101101111110111011110101001110101011;
          9:
            level_vec_out = 64'b0111011111011111000001110111101101111110111011110101001110101011;
          10:
            level_vec_out = 64'b0111011111011111000001110111101101111110111011110101001110111011;
          11:
            level_vec_out = 64'b0111011111011111000001110111101101111110111011110101011110111011;
          12:
            level_vec_out = 64'b0111011111011111010001110111101101111110111011110101011110111011;
          13:
            level_vec_out = 64'b0111011111011111010001110111101101111110111011110101011111111011;
          14:
            level_vec_out = 64'b0111011111011111010001110111101101111110111011110101011111111011;
          15:
            level_vec_out = 64'b0111011111011111010001110111101101111110111011110101011111111011;
          16:
            level_vec_out = 64'b1111011111011111010001110111101101111110111011110101011111111011;
          17:
            level_vec_out = 64'b1111011111011111010001110111101101111110111011110101111111111011;
          18:
            level_vec_out = 64'b1111011111011111010001110111101101111110111011110101111111111011;
          19:
            level_vec_out = 64'b1111011111011111010001110111101101111110111011110101111111111011;
          20:
            level_vec_out = 64'b1111011111011111011001110111101101111110111011110101111111111011;
          21:
            level_vec_out = 64'b1111011111111111011001110111101101111110111011110101111111111011;
          22:
            level_vec_out = 64'b1111011111111111011101110111101101111110111011110101111111111011;
          23:
            level_vec_out = 64'b1111111111111111011101111111101101111110111011110101111111111111;
          24:
            level_vec_out = 64'b1111111111111111011101111111101111111110111011111101111111111111;
          25:
            level_vec_out = 64'b1111111111111111011101111111111111111111111111111101111111111111;
          26:
            level_vec_out = 64'b1111111111111111011101111111111111111111111111111101111111111111;
          27:
            level_vec_out = 64'b1111111111111111011101111111111111111111111111111101111111111111;
          28:
            level_vec_out = 64'b1111111111111111011101111111111111111111111111111101111111111111;
          29:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111101111111111111;
          30:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111101111111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111101111111111111;
        endcase
      6:
        case (frame_id)
          0:
            level_vec_out = 64'b1111011001001111011100001111010001011101011111000100110010010110;
          1:
            level_vec_out = 64'b1111011001001111011100001111010001011101011111000100110010010110;
          2:
            level_vec_out = 64'b1111011001001111011101001111010001011101011111000100110010110110;
          3:
            level_vec_out = 64'b1111011001001111011101001111010001011101011111000100110010110110;
          4:
            level_vec_out = 64'b1111011011001111011101001111010011011101011111010100111010110110;
          5:
            level_vec_out = 64'b1111011011001111011101001111010011011101011111010100111010110110;
          6:
            level_vec_out = 64'b1111011011001111011111001111010011011101011111010100111010110110;
          7:
            level_vec_out = 64'b1111011011001111011111001111010011111101011111010100111010110110;
          8:
            level_vec_out = 64'b1111011011001111011111001111010011111101011111010101111010110110;
          9:
            level_vec_out = 64'b1111011011101111011111001111110011111101011111010101111010110110;
          10:
            level_vec_out = 64'b1111011011101111011111001111110011111101011111010111111010110110;
          11:
            level_vec_out = 64'b1111011011101111111111011111111111111101011111010111111010110110;
          12:
            level_vec_out = 64'b1111011011101111111111011111111111111101011111010111111010110110;
          13:
            level_vec_out = 64'b1111011011111111111111011111111111111101011111010111111010110110;
          14:
            level_vec_out = 64'b1111011011111111111111011111111111111101011111010111111010110110;
          15:
            level_vec_out = 64'b1111011011111111111111011111111111111101011111010111111010110110;
          16:
            level_vec_out = 64'b1111011011111111111111011111111111111101011111010111111010111110;
          17:
            level_vec_out = 64'b1111011011111111111111011111111111111101111111010111111010111110;
          18:
            level_vec_out = 64'b1111111011111111111111011111111111111101111111010111111010111110;
          19:
            level_vec_out = 64'b1111111011111111111111011111111111111101111111010111111010111110;
          20:
            level_vec_out = 64'b1111111011111111111111011111111111111101111111010111111010111110;
          21:
            level_vec_out = 64'b1111111011111111111111111111111111111101111111010111111010111110;
          22:
            level_vec_out = 64'b1111111011111111111111111111111111111111111111010111111010111110;
          23:
            level_vec_out = 64'b1111111011111111111111111111111111111111111111010111111011111110;
          24:
            level_vec_out = 64'b1111111011111111111111111111111111111111111111010111111011111110;
          25:
            level_vec_out = 64'b1111111011111111111111111111111111111111111111010111111111111110;
          26:
            level_vec_out = 64'b1111111011111111111111111111111111111111111111010111111111111110;
          27:
            level_vec_out = 64'b1111111011111111111111111111111111111111111111010111111111111111;
          28:
            level_vec_out = 64'b1111111011111111111111111111111111111111111111010111111111111111;
          29:
            level_vec_out = 64'b1111111011111111111111111111111111111111111111010111111111111111;
          30:
            level_vec_out = 64'b1111111011111111111111111111111111111111111111111111111111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        endcase
      7:
        case (frame_id)
          0:
            level_vec_out = 64'b0011110001010011100011001100100001000111000110000001000000101111;
          1:
            level_vec_out = 64'b0011110001011011100011001100100001100111000110000001000000101111;
          2:
            level_vec_out = 64'b0011110001011011100011001100100001100111000110000001000000101111;
          3:
            level_vec_out = 64'b0011110001011011100011001110100001101111000110000001000000101111;
          4:
            level_vec_out = 64'b0011110001111011110011001110100001101111000110000101000000101111;
          5:
            level_vec_out = 64'b0011110001111011110011001110100001101111000110000101000000101111;
          6:
            level_vec_out = 64'b0011110001111011110011001110100001101111000110000101000000101111;
          7:
            level_vec_out = 64'b0011110001111011110011001110100001101111000111010101000000101111;
          8:
            level_vec_out = 64'b0011110001111011110011001110100001101111000111010101000000101111;
          9:
            level_vec_out = 64'b0111110101111011110011001110100001101111000111010101000000101111;
          10:
            level_vec_out = 64'b0111110101111011110011001110100011101111000111010101000100101111;
          11:
            level_vec_out = 64'b0111110101111011110011101110100011101111000111010101000110101111;
          12:
            level_vec_out = 64'b0111110101111011111011111110100011101111000111010101000110101111;
          13:
            level_vec_out = 64'b0111110101111011111011111110100011101111000111010101000110101111;
          14:
            level_vec_out = 64'b0111110101111011111011111110100011101111000111010101000110101111;
          15:
            level_vec_out = 64'b0111110101111011111011111110100011101111000111010101000110101111;
          16:
            level_vec_out = 64'b0111110101111011111011111110101011101111100111010101000110101111;
          17:
            level_vec_out = 64'b0111110101111011111011111110101011101111100111010101000110101111;
          18:
            level_vec_out = 64'b0111111101111011111011111110101011101111100111110101000110101111;
          19:
            level_vec_out = 64'b0111111101111011111011111110101011101111100111110101000110101111;
          20:
            level_vec_out = 64'b0111111101111111111011111110101011101111100111110101000110101111;
          21:
            level_vec_out = 64'b0111111101111111111011111110101011101111100111110101000110111111;
          22:
            level_vec_out = 64'b0111111101111111111011111110101011101111100111110101000110111111;
          23:
            level_vec_out = 64'b1111111101111111111011111110101011101111100111110101010110111111;
          24:
            level_vec_out = 64'b1111111111111111111011111110111011101111100111110101010110111111;
          25:
            level_vec_out = 64'b1111111111111111111011111110111011101111100111110101010110111111;
          26:
            level_vec_out = 64'b1111111111111111111011111110111011101111101111110101011110111111;
          27:
            level_vec_out = 64'b1111111111111111111011111111111011111111101111111101011110111111;
          28:
            level_vec_out = 64'b1111111111111111111011111111111111111111101111111111111110111111;
          29:
            level_vec_out = 64'b1111111111111111111011111111111111111111101111111111111110111111;
          30:
            level_vec_out = 64'b1111111111111111111011111111111111111111101111111111111110111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        endcase
    endcase
  end
endmodule