/**
 * @file level_hvec_gen_hdl.hpp
 * @brief This script generates HDL code for generating high-dimensional LEVEL vectors.
 * It is a novel method; for more information, please refer to our paper.
 *
 * @author Saeid Jamili and Marco Angioli
 * @note Author names are listed in alphabetical order.
 * @email <saeid.jamili@uniroma1.it>
 * @email <marco.angioli@uniroma1.it>
 *
 * @contributors
 *
 * @date Created: 24th July 2023
 * @date Last Updated: 23th August 2023
 *
 * @version 1.0.0
 *
 * @institute Sapienza University of Rome
 * @cite https://doi.org/10.xxxx/yyyyy
 *
 * @section DEPENDENCIES
 * - Dependency1: Description or version details.
 * - Dependency2: Description or version details.
 *
 * @section LICENSE
 * This file is part of the Aeneas HyperCompute Platform.
 *
 * Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 *
 * @section CHANGELOG
 * @version 1.0.0-dev - 23th August 2023
 * - Initial release
 *
 * @todo
 * - Complete level vector generator function
 * - Add training
 *
 * @see
 * -
 * -
 * -
 *
 */

module level_hvec_gen #(parameter int DI_PARALLEL_W_BITS = 64) (
  input logic [2:0] frame_index,
  input logic [4:0] frame_id,
  output logic [DI_PARALLEL_W_BITS-1:0] level_vec_out
);
  always_comb begin
    case (frame_index)
      0:
        case (frame_id)
          0:
            level_vec_out = 64'b0010010110001110001011101111110000101111010011101100010110001010;
          1:
            level_vec_out = 64'b0010010110001110001011101111110000101111010011101100010110001010;
          2:
            level_vec_out = 64'b0010110110001110001011101111110000101111010011101100010110001010;
          3:
            level_vec_out = 64'b0010110111001110001011101111110000101111010011101100010110001010;
          4:
            level_vec_out = 64'b0010110111001110001011101111110000101111010011101100010110001010;
          5:
            level_vec_out = 64'b0010110111001110001011101111110000111111010011101100010110001010;
          6:
            level_vec_out = 64'b1110110111001110001011101111110000111111011011101100010110001010;
          7:
            level_vec_out = 64'b1110110111001110001011101111110000111111011011101100010110001010;
          8:
            level_vec_out = 64'b1110110111001110001011101111111000111111011011101100010110001110;
          9:
            level_vec_out = 64'b1110110111001110001011101111111000111111011011101100010111001110;
          10:
            level_vec_out = 64'b1110110111001110001011101111111000111111011011101100110111001110;
          11:
            level_vec_out = 64'b1110110111001110001011101111111000111111011011101100110111001111;
          12:
            level_vec_out = 64'b1110110111001110001011111111111000111111011011101100110111001111;
          13:
            level_vec_out = 64'b1110110111001110001011111111111000111111011011101110110111001111;
          14:
            level_vec_out = 64'b1110110111001110001011111111111000111111011011101110110111011111;
          15:
            level_vec_out = 64'b1110110111001110101011111111111000111111011011101110110111011111;
          16:
            level_vec_out = 64'b1110110111101110101011111111111000111111011011101110110111111111;
          17:
            level_vec_out = 64'b1110110111101110101011111111111010111111011111101110110111111111;
          18:
            level_vec_out = 64'b1110110111101110101011111111111010111111011111111110111111111111;
          19:
            level_vec_out = 64'b1110110111101110101011111111111010111111011111111110111111111111;
          20:
            level_vec_out = 64'b1110110111101110101011111111111010111111011111111110111111111111;
          21:
            level_vec_out = 64'b1110110111101110101011111111111010111111011111111110111111111111;
          22:
            level_vec_out = 64'b1110110111101110101011111111111010111111111111111111111111111111;
          23:
            level_vec_out = 64'b1110110111101111101011111111111010111111111111111111111111111111;
          24:
            level_vec_out = 64'b1110110111101111101011111111111011111111111111111111111111111111;
          25:
            level_vec_out = 64'b1110110111101111101011111111111011111111111111111111111111111111;
          26:
            level_vec_out = 64'b1110111111111111101011111111111011111111111111111111111111111111;
          27:
            level_vec_out = 64'b1110111111111111101011111111111011111111111111111111111111111111;
          28:
            level_vec_out = 64'b1110111111111111101111111111111011111111111111111111111111111111;
          29:
            level_vec_out = 64'b1111111111111111101111111111111011111111111111111111111111111111;
          30:
            level_vec_out = 64'b1111111111111111101111111111111111111111111111111111111111111111;
          31:
            level_vec_out = 64'b1111111111111111101111111111111111111111111111111111111111111111;
        endcase
      1:
        case (frame_id)
          0:
            level_vec_out = 64'b0011100000010100100000100011100100011110001101110001111111111100;
          1:
            level_vec_out = 64'b0011100000010100100000100011100100011110001101110001111111111101;
          2:
            level_vec_out = 64'b0011100000010100100010100011100100011110011101110001111111111101;
          3:
            level_vec_out = 64'b0011100001010100100010100011100100011110011101110001111111111101;
          4:
            level_vec_out = 64'b0011100001010110100110100011100100011110011101110001111111111101;
          5:
            level_vec_out = 64'b0011100001110110100110100011100100011110011101110001111111111101;
          6:
            level_vec_out = 64'b0011100001110110100110100011100100011110011101110001111111111101;
          7:
            level_vec_out = 64'b0011100001110110100110100011100100011110011101110001111111111101;
          8:
            level_vec_out = 64'b0011100001110110100110100011100100011110011101110001111111111101;
          9:
            level_vec_out = 64'b0011100001110110100110100011110100011110011111110001111111111101;
          10:
            level_vec_out = 64'b0011100001110110100110101011111100011110011111110001111111111101;
          11:
            level_vec_out = 64'b0011101001110110100110101011111100011110011111110001111111111101;
          12:
            level_vec_out = 64'b0011101001110110100110101011111100111110011111110001111111111101;
          13:
            level_vec_out = 64'b0011101001110110100110101011111100111110011111110001111111111101;
          14:
            level_vec_out = 64'b0011101001110110100110101011111100111110111111110001111111111101;
          15:
            level_vec_out = 64'b0011101001110110100110101011111101111110111111110001111111111101;
          16:
            level_vec_out = 64'b0011101001110110100110101011111101111110111111110001111111111101;
          17:
            level_vec_out = 64'b0011101001110110100110101111111101111110111111110001111111111101;
          18:
            level_vec_out = 64'b0011101011111110100110111111111101111110111111110011111111111101;
          19:
            level_vec_out = 64'b0111101011111110100110111111111101111111111111111011111111111101;
          20:
            level_vec_out = 64'b0111101011111110100110111111111101111111111111111011111111111101;
          21:
            level_vec_out = 64'b0111101111111110100110111111111101111111111111111011111111111101;
          22:
            level_vec_out = 64'b0111101111111110100110111111111101111111111111111011111111111101;
          23:
            level_vec_out = 64'b0111101111111110100110111111111101111111111111111011111111111101;
          24:
            level_vec_out = 64'b0111101111111110100110111111111101111111111111111011111111111101;
          25:
            level_vec_out = 64'b0111101111111110110110111111111101111111111111111011111111111101;
          26:
            level_vec_out = 64'b1111101111111110110110111111111101111111111111111011111111111101;
          27:
            level_vec_out = 64'b1111101111111111110110111111111101111111111111111011111111111101;
          28:
            level_vec_out = 64'b1111101111111111110111111111111111111111111111111011111111111101;
          29:
            level_vec_out = 64'b1111101111111111110111111111111111111111111111111111111111111101;
          30:
            level_vec_out = 64'b1111111111111111110111111111111111111111111111111111111111111101;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111101;
        endcase
      2:
        case (frame_id)
          0:
            level_vec_out = 64'b1001111111110010110001101100111110110000011010111101010110111110;
          1:
            level_vec_out = 64'b1001111111110010110001101100111110110000011010111101010110111110;
          2:
            level_vec_out = 64'b1001111111110010110001101100111110110000011010111101010110111110;
          3:
            level_vec_out = 64'b1001111111110010110001101100111110110010011010111101010110111110;
          4:
            level_vec_out = 64'b1001111111110010110001111100111110110010011010111101010110111110;
          5:
            level_vec_out = 64'b1001111111110010110001111100111110110010011010111101010110111110;
          6:
            level_vec_out = 64'b1001111111110010110001111100111111110010011010111101010110111110;
          7:
            level_vec_out = 64'b1001111111110010110001111100111111110010111010111101010110111110;
          8:
            level_vec_out = 64'b1001111111110010111001111100111111110010111010111101010110111110;
          9:
            level_vec_out = 64'b1001111111110010111001111110111111110010111010111101010110111110;
          10:
            level_vec_out = 64'b1001111111110010111001111110111111110010111010111101010110111110;
          11:
            level_vec_out = 64'b1001111111110010111001111110111111110010111010111111010110111110;
          12:
            level_vec_out = 64'b1001111111110010111101111110111111110010111010111111010110111110;
          13:
            level_vec_out = 64'b1001111111110010111101111110111111110010111110111111010110111110;
          14:
            level_vec_out = 64'b1101111111110010111101111110111111111010111110111111011110111110;
          15:
            level_vec_out = 64'b1101111111110010111101111110111111111010111110111111011111111111;
          16:
            level_vec_out = 64'b1101111111110010111101111110111111111010111110111111011111111111;
          17:
            level_vec_out = 64'b1101111111110010111101111110111111111010111111111111011111111111;
          18:
            level_vec_out = 64'b1101111111110010111101111110111111111010111111111111011111111111;
          19:
            level_vec_out = 64'b1101111111110011111101111110111111111010111111111111011111111111;
          20:
            level_vec_out = 64'b1101111111110011111101111111111111111010111111111111011111111111;
          21:
            level_vec_out = 64'b1101111111110011111101111111111111111010111111111111011111111111;
          22:
            level_vec_out = 64'b1101111111110011111101111111111111111010111111111111011111111111;
          23:
            level_vec_out = 64'b1101111111110111111101111111111111111010111111111111011111111111;
          24:
            level_vec_out = 64'b1101111111110111111101111111111111111010111111111111011111111111;
          25:
            level_vec_out = 64'b1101111111110111111101111111111111111110111111111111011111111111;
          26:
            level_vec_out = 64'b1101111111110111111111111111111111111110111111111111011111111111;
          27:
            level_vec_out = 64'b1101111111110111111111111111111111111110111111111111011111111111;
          28:
            level_vec_out = 64'b1101111111110111111111111111111111111110111111111111011111111111;
          29:
            level_vec_out = 64'b1101111111111111111111111111111111111110111111111111011111111111;
          30:
            level_vec_out = 64'b1101111111111111111111111111111111111110111111111111011111111111;
          31:
            level_vec_out = 64'b1101111111111111111111111111111111111111111111111111011111111111;
        endcase
      3:
        case (frame_id)
          0:
            level_vec_out = 64'b1001100011001001010000100101101001100011010100100111100110000001;
          1:
            level_vec_out = 64'b1001100011001001010100100101101001100111010100100111101110001001;
          2:
            level_vec_out = 64'b1001100011001001110100100101101001100111010100100111101110001001;
          3:
            level_vec_out = 64'b1001100011001101110100100101101001100111010100100111101110001001;
          4:
            level_vec_out = 64'b1001100011001101110100100101111001100111010100100111111110001001;
          5:
            level_vec_out = 64'b1001100011001101110100100101111101100111010101100111111110001001;
          6:
            level_vec_out = 64'b1001100111001101110100100101111101100111010101100111111110001001;
          7:
            level_vec_out = 64'b1001100111101101110100100101111101100111010101100111111110001001;
          8:
            level_vec_out = 64'b1001100111101101110100100101111101100111010101100111111110001001;
          9:
            level_vec_out = 64'b1001100111101101111100100111111101100111010101100111111110001001;
          10:
            level_vec_out = 64'b1001100111101101111100100111111101100111010101100111111110001001;
          11:
            level_vec_out = 64'b1001100111101101111100100111111101100111110101100111111110001001;
          12:
            level_vec_out = 64'b1101100111101101111100100111111101100111110101100111111110001001;
          13:
            level_vec_out = 64'b1101100111101101111110100111111101100111110101110111111110101001;
          14:
            level_vec_out = 64'b1101100111101101111110100111111101100111110101110111111110101001;
          15:
            level_vec_out = 64'b1101101111101101111110100111111101100111110101110111111110101001;
          16:
            level_vec_out = 64'b1101101111101101111110100111111101100111110101110111111110101101;
          17:
            level_vec_out = 64'b1101101111101101111110100111111101100111110101110111111110101101;
          18:
            level_vec_out = 64'b1101101111101101111110100111111101100111110101110111111110101101;
          19:
            level_vec_out = 64'b1101101111101101111110110111111101100111110101110111111110101101;
          20:
            level_vec_out = 64'b1101101111101101111110110111111101100111110101110111111110111101;
          21:
            level_vec_out = 64'b1101111111101101111110110111111101100111110101110111111110111101;
          22:
            level_vec_out = 64'b1101111111101101111110110111111101100111110101110111111110111101;
          23:
            level_vec_out = 64'b1101111111101101111110110111111101100111111101110111111111111101;
          24:
            level_vec_out = 64'b1101111111101111111110110111111101100111111101111111111111111111;
          25:
            level_vec_out = 64'b1101111111101111111110111111111101100111111101111111111111111111;
          26:
            level_vec_out = 64'b1101111111101111111110111111111101100111111101111111111111111111;
          27:
            level_vec_out = 64'b1101111111101111111110111111111101110111111111111111111111111111;
          28:
            level_vec_out = 64'b1101111111111111111111111111111101111111111111111111111111111111;
          29:
            level_vec_out = 64'b1101111111111111111111111111111111111111111111111111111111111111;
          30:
            level_vec_out = 64'b1101111111111111111111111111111111111111111111111111111111111111;
          31:
            level_vec_out = 64'b1101111111111111111111111111111111111111111111111111111111111111;
        endcase
      4:
        case (frame_id)
          0:
            level_vec_out = 64'b0001011110101100001111000100111001110101011111001111101101011011;
          1:
            level_vec_out = 64'b0001011110101100001111000100111001110101011111001111101101011111;
          2:
            level_vec_out = 64'b0001011110101100001111000100111011110101011111001111101101011111;
          3:
            level_vec_out = 64'b0001011110101100001111000100111011110101011111001111101101011111;
          4:
            level_vec_out = 64'b0001011110101100001111000100111011110111011111001111101101011111;
          5:
            level_vec_out = 64'b0001011110101101001111000100111011110111111111001111101101011111;
          6:
            level_vec_out = 64'b0001011110101101001111000110111011110111111111001111101101011111;
          7:
            level_vec_out = 64'b0001011110101101001111000110111011110111111111001111101101011111;
          8:
            level_vec_out = 64'b0001011110101101001111000110111011110111111111001111101101011111;
          9:
            level_vec_out = 64'b0001011110101101001111000110111011110111111111001111101101011111;
          10:
            level_vec_out = 64'b0001011111101101001111000110111111110111111111001111101101011111;
          11:
            level_vec_out = 64'b0001011111101101001111000110111111110111111111001111101101011111;
          12:
            level_vec_out = 64'b0001011111101101001111000110111111110111111111001111101101011111;
          13:
            level_vec_out = 64'b0001011111101101001111000110111111110111111111001111101101011111;
          14:
            level_vec_out = 64'b0001011111101101001111000110111111110111111111001111101101011111;
          15:
            level_vec_out = 64'b0011011111101101001111000110111111110111111111001111101101011111;
          16:
            level_vec_out = 64'b0011011111101101001111000110111111110111111111001111101101011111;
          17:
            level_vec_out = 64'b0011011111101101001111100111111111110111111111001111101101011111;
          18:
            level_vec_out = 64'b0011011111101101001111100111111111110111111111001111101101011111;
          19:
            level_vec_out = 64'b0011011111101101001111100111111111110111111111001111101101011111;
          20:
            level_vec_out = 64'b0011011111101101001111100111111111110111111111001111111101011111;
          21:
            level_vec_out = 64'b0011011111101101001111100111111111110111111111001111111101011111;
          22:
            level_vec_out = 64'b0011011111101101111111100111111111110111111111001111111101011111;
          23:
            level_vec_out = 64'b0011011111101101111111100111111111110111111111001111111101111111;
          24:
            level_vec_out = 64'b0011011111101101111111100111111111110111111111001111111101111111;
          25:
            level_vec_out = 64'b0011011111101101111111100111111111110111111111101111111101111111;
          26:
            level_vec_out = 64'b0011011111111101111111110111111111110111111111101111111101111111;
          27:
            level_vec_out = 64'b1111011111111111111111110111111111110111111111101111111101111111;
          28:
            level_vec_out = 64'b1111011111111111111111110111111111111111111111101111111101111111;
          29:
            level_vec_out = 64'b1111011111111111111111110111111111111111111111101111111101111111;
          30:
            level_vec_out = 64'b1111011111111111111111111111111111111111111111101111111111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        endcase
      5:
        case (frame_id)
          0:
            level_vec_out = 64'b0101101001100110100110000010011001011111011110110100110101001100;
          1:
            level_vec_out = 64'b0101101001110110100110000010011001011111011110110100110101001100;
          2:
            level_vec_out = 64'b0101101001110110100110000010011101011111011110110100110101001100;
          3:
            level_vec_out = 64'b0101101001110110100110000010011101011111011110110100110101001100;
          4:
            level_vec_out = 64'b0101101001110110100110000010011101011111011110110100110101001100;
          5:
            level_vec_out = 64'b0101111001110110100110000010011101011111011110110100110101001100;
          6:
            level_vec_out = 64'b0101111001110110100110000010011101011111011110110100110101001100;
          7:
            level_vec_out = 64'b0101111001110110110110001010011101011111011110110100110101001100;
          8:
            level_vec_out = 64'b0111111001110110110110001011011101011111011110110100110101101100;
          9:
            level_vec_out = 64'b1111111001110110110110001011011101011111011110110100110101101100;
          10:
            level_vec_out = 64'b1111111001110110110110011011011101011111011110110100110101101110;
          11:
            level_vec_out = 64'b1111111001110110110110111011011101011111011110110100110111101110;
          12:
            level_vec_out = 64'b1111111001110110110110111011011101011111011110110101110111101110;
          13:
            level_vec_out = 64'b1111111001110110110110111111011101011111011110110101110111101110;
          14:
            level_vec_out = 64'b1111111001110110110110111111011111011111011110110101110111111110;
          15:
            level_vec_out = 64'b1111111001110110110110111111011111011111011110110101110111111110;
          16:
            level_vec_out = 64'b1111111001110110110110111111011111011111011110111101110111111110;
          17:
            level_vec_out = 64'b1111111001110110110111111111011111011111011110111101110111111110;
          18:
            level_vec_out = 64'b1111111001110110110111111111011111011111011110111101110111111110;
          19:
            level_vec_out = 64'b1111111001110110110111111111011111111111011110111111110111111110;
          20:
            level_vec_out = 64'b1111111101110110110111111111111111111111011110111111110111111110;
          21:
            level_vec_out = 64'b1111111111110110110111111111111111111111011110111111110111111110;
          22:
            level_vec_out = 64'b1111111111110110110111111111111111111111011110111111110111111110;
          23:
            level_vec_out = 64'b1111111111110110110111111111111111111111011110111111110111111110;
          24:
            level_vec_out = 64'b1111111111110110110111111111111111111111011110111111111111111110;
          25:
            level_vec_out = 64'b1111111111110110110111111111111111111111011111111111111111111110;
          26:
            level_vec_out = 64'b1111111111110111110111111111111111111111011111111111111111111110;
          27:
            level_vec_out = 64'b1111111111111111111111111111111111111111011111111111111111111110;
          28:
            level_vec_out = 64'b1111111111111111111111111111111111111111011111111111111111111110;
          29:
            level_vec_out = 64'b1111111111111111111111111111111111111111011111111111111111111110;
          30:
            level_vec_out = 64'b1111111111111111111111111111111111111111011111111111111111111110;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111011111111111111111111111;
        endcase
      6:
        case (frame_id)
          0:
            level_vec_out = 64'b1101010000000111000100110011110000100010111100000100111001101100;
          1:
            level_vec_out = 64'b1101010000000111000100110011110000100010111100000100111001101100;
          2:
            level_vec_out = 64'b1101010000000111000100110111110000100110111100000100111001101100;
          3:
            level_vec_out = 64'b1101010100000111000100110111110000100110111100000100111101101100;
          4:
            level_vec_out = 64'b1101010100000111000100110111110000100110111100000110111111101100;
          5:
            level_vec_out = 64'b1101010100000111000100110111110000100110111100000110111111101100;
          6:
            level_vec_out = 64'b1101010110000111000100110111110000100110111100000110111111101100;
          7:
            level_vec_out = 64'b1111010110000111000100110111110000100110111100000110111111101100;
          8:
            level_vec_out = 64'b1111010110000111000100110111110000100110111100000110111111101101;
          9:
            level_vec_out = 64'b1111010110000111000100110111110000100110111110000110111111101101;
          10:
            level_vec_out = 64'b1111010110000111000101110111110000100110111110000110111111101101;
          11:
            level_vec_out = 64'b1111010110000111000101110111110100100110111110000110111111101101;
          12:
            level_vec_out = 64'b1111010110001111000101110111110101100110111110000110111111101101;
          13:
            level_vec_out = 64'b1111010110011111000101110111110101101110111110000110111111101101;
          14:
            level_vec_out = 64'b1111010110011111000101110111110101101110111110000110111111101101;
          15:
            level_vec_out = 64'b1111010110011111000101110111110101101110111110001110111111101101;
          16:
            level_vec_out = 64'b1111010110011111000101110111110101101110111110001110111111101101;
          17:
            level_vec_out = 64'b1111010110011111000101110111110101101110111111001110111111101101;
          18:
            level_vec_out = 64'b1111010110011111000101110111111101101110111111001110111111101111;
          19:
            level_vec_out = 64'b1111010111011111000101110111111101101110111111001110111111101111;
          20:
            level_vec_out = 64'b1111010111011111000101110111111101101110111111001110111111101111;
          21:
            level_vec_out = 64'b1111110111011111000101110111111101111110111111001110111111101111;
          22:
            level_vec_out = 64'b1111110111011111000101111111111111111110111111001110111111101111;
          23:
            level_vec_out = 64'b1111110111011111100101111111111111111110111111001111111111101111;
          24:
            level_vec_out = 64'b1111110111011111100111111111111111111110111111001111111111101111;
          25:
            level_vec_out = 64'b1111110111011111110111111111111111111110111111011111111111101111;
          26:
            level_vec_out = 64'b1111110111011111111111111111111111111110111111011111111111101111;
          27:
            level_vec_out = 64'b1111110111011111111111111111111111111110111111011111111111101111;
          28:
            level_vec_out = 64'b1111111111011111111111111111111111111110111111011111111111101111;
          29:
            level_vec_out = 64'b1111111111011111111111111111111111111110111111011111111111101111;
          30:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111011111111111101111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111011111111111111111;
        endcase
      7:
        case (frame_id)
          0:
            level_vec_out = 64'b1001110100000101000100110110101000010000000110011011100000101101;
          1:
            level_vec_out = 64'b1001110100000101000100110110101010010000000110011011100000101101;
          2:
            level_vec_out = 64'b1001110100000101000100110110101010010000000110011011100000101101;
          3:
            level_vec_out = 64'b1101111100000101000100110110101010010000000110011011100000101101;
          4:
            level_vec_out = 64'b1101111100000101000100110110101010010000000110011011100000101101;
          5:
            level_vec_out = 64'b1101111100000101000100110110101010010000000110011111100000101101;
          6:
            level_vec_out = 64'b1101111100000101000100110110101010010000000110011111100000101111;
          7:
            level_vec_out = 64'b1101111100000101000100111110101110010000000110011111100001101111;
          8:
            level_vec_out = 64'b1101111100000101000100111110101110010000100110011111100001101111;
          9:
            level_vec_out = 64'b1101111100000101000100111110101110010000100110011111100001101111;
          10:
            level_vec_out = 64'b1101111100000101000100111110101110010000100110011111100001101111;
          11:
            level_vec_out = 64'b1101111100000101000100111110101110010000100110011111101001101111;
          12:
            level_vec_out = 64'b1111111100000101000100111110101110010000100110011111101001101111;
          13:
            level_vec_out = 64'b1111111100000101000100111110101110010000100110011111101001101111;
          14:
            level_vec_out = 64'b1111111100000101000100111110101110010000100111011111101001101111;
          15:
            level_vec_out = 64'b1111111100000101000100111110101111010000100111011111101001101111;
          16:
            level_vec_out = 64'b1111111100010101000100111111101111010010101111011111101001101111;
          17:
            level_vec_out = 64'b1111111100010101000100111111101111010010101111011111101001101111;
          18:
            level_vec_out = 64'b1111111100010101000100111111101111010010101111011111101001101111;
          19:
            level_vec_out = 64'b1111111100010101000100111111101111010010101111011111101001101111;
          20:
            level_vec_out = 64'b1111111110010101000100111111101111010010101111111111101001111111;
          21:
            level_vec_out = 64'b1111111110010101010101111111111111010010101111111111101001111111;
          22:
            level_vec_out = 64'b1111111111010101010101111111111111010011101111111111101001111111;
          23:
            level_vec_out = 64'b1111111111010101010101111111111111110011101111111111101001111111;
          24:
            level_vec_out = 64'b1111111111010101011101111111111111111011101111111111101001111111;
          25:
            level_vec_out = 64'b1111111111010101011101111111111111111011101111111111101011111111;
          26:
            level_vec_out = 64'b1111111111010101011101111111111111111011101111111111101011111111;
          27:
            level_vec_out = 64'b1111111111010101011101111111111111111011101111111111101011111111;
          28:
            level_vec_out = 64'b1111111111010101011101111111111111111011101111111111101011111111;
          29:
            level_vec_out = 64'b1111111111010101111101111111111111111111111111111111111011111111;
          30:
            level_vec_out = 64'b1111111111111101111101111111111111111111111111111111111011111111;
          31:
            level_vec_out = 64'b1111111111111101111111111111111111111111111111111111111111111111;
        endcase
    endcase
  end
endmodule