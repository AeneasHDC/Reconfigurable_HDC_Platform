/**
 * @file level_hvec_gen_hdl.hpp
 * @brief This script generates HDL code for generating high-dimensional LEVEL vectors.
 * It is a novel method; for more information, please refer to our paper.
 *
 * @author Saeid Jamili and Marco Angioli
 * @note Author names are listed in alphabetical order.
 * @email <saeid.jamili@uniroma1.it>
 * @email <marco.angioli@uniroma1.it>
 *
 * @contributors
 *
 * @date Created: 24th July 2023
 * @date Last Updated: 23th August 2023
 *
 * @version 1.0.0
 *
 * @institute Sapienza University of Rome
 * @cite https://doi.org/10.xxxx/yyyyy
 *
 * @section DEPENDENCIES
 * - Dependency1: Description or version details.
 * - Dependency2: Description or version details.
 *
 * @section LICENSE
 * This file is part of the Aeneas HyperCompute Platform.
 *
 * Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 *
 * @section CHANGELOG
 * @version 1.0.0-dev - 23th August 2023
 * - Initial release
 *
 * @todo
 * - Complete level vector generator function
 * - Add training
 *
 * @see
 * -
 * -
 * -
 *
 */

module level_hvec_gen #(parameter int DI_PARALLEL_W_BITS = 64) (
  input logic [2:0] frame_index,
  input logic [4:0] frame_id,
  output logic [DI_PARALLEL_W_BITS-1:0] level_vec_out
);
  always_comb begin
    case (frame_index)
      0:
        case (frame_id)
          0:
            level_vec_out = 64'b0000110101011001011101011011100100010001111010101101000100100000;
          1:
            level_vec_out = 64'b1000110101011001011101111011100100010001111010101101000100100000;
          2:
            level_vec_out = 64'b1000111101011001011101111011100100010001111010111101000100100000;
          3:
            level_vec_out = 64'b1000111101011001011101111011100100010001111010111101000100100010;
          4:
            level_vec_out = 64'b1000111101011011011111111011100100010001111010111101000100100010;
          5:
            level_vec_out = 64'b1000111101011011011111111011110100010001111010111101000100100010;
          6:
            level_vec_out = 64'b1000111101011011011111111011110100010001111110111111000100100010;
          7:
            level_vec_out = 64'b1000111101011011011111111011110101011001111110111111000100100010;
          8:
            level_vec_out = 64'b1000111101011011011111111011110101011001111110111111000100100010;
          9:
            level_vec_out = 64'b1000111101011011011111111011110101011001111110111111000100100010;
          10:
            level_vec_out = 64'b1000111101011011011111111011110101011001111110111111000100100010;
          11:
            level_vec_out = 64'b1000111101011011011111111011110101011001111110111111000100100010;
          12:
            level_vec_out = 64'b1000111101011011011111111011110101011001111110111111000100100010;
          13:
            level_vec_out = 64'b1001111101011011011111111011110101011001111110111111000100100010;
          14:
            level_vec_out = 64'b1001111101011011111111111011110101011001111110111111000100100010;
          15:
            level_vec_out = 64'b1001111101011011111111111011111101011101111110111111000100100010;
          16:
            level_vec_out = 64'b1001111101011011111111111011111101011101111110111111000110100010;
          17:
            level_vec_out = 64'b1001111101011011111111111011111101011101111111111111000110110010;
          18:
            level_vec_out = 64'b1001111101011011111111111011111101011101111111111111000110110010;
          19:
            level_vec_out = 64'b1001111111011011111111111011111101011101111111111111000110110010;
          20:
            level_vec_out = 64'b1011111111011011111111111011111111011101111111111111000110110010;
          21:
            level_vec_out = 64'b1011111111111011111111111111111111011101111111111111001110110010;
          22:
            level_vec_out = 64'b1011111111111011111111111111111111011101111111111111001110110010;
          23:
            level_vec_out = 64'b1111111111111011111111111111111111011101111111111111001111110010;
          24:
            level_vec_out = 64'b1111111111111011111111111111111111111101111111111111001111110010;
          25:
            level_vec_out = 64'b1111111111111011111111111111111111111101111111111111001111110011;
          26:
            level_vec_out = 64'b1111111111111011111111111111111111111111111111111111001111110011;
          27:
            level_vec_out = 64'b1111111111111011111111111111111111111111111111111111011111110011;
          28:
            level_vec_out = 64'b1111111111111011111111111111111111111111111111111111011111110011;
          29:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111011111110011;
          30:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111011111110111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        endcase
      1:
        case (frame_id)
          0:
            level_vec_out = 64'b0110001110010010100111110111010100110001011110111101110110011001;
          1:
            level_vec_out = 64'b1110001110010111100111110111010100110001011110111101110110011001;
          2:
            level_vec_out = 64'b1110001110010111100111110111010100110001011110111101110110011001;
          3:
            level_vec_out = 64'b1110001110010111100111110111010100110001111110111101110110011001;
          4:
            level_vec_out = 64'b1110001111010111100111110111010110110001111110111101110110011001;
          5:
            level_vec_out = 64'b1110001111010111100111110111010110110001111110111101110110011001;
          6:
            level_vec_out = 64'b1110001111010111100111110111010110111101111110111101110110011001;
          7:
            level_vec_out = 64'b1110001111010111110111110111010110111101111110111101110110011001;
          8:
            level_vec_out = 64'b1110001111010111110111110111010110111101111110111101110110011001;
          9:
            level_vec_out = 64'b1110001111010111110111110111010110111101111110111101110110011001;
          10:
            level_vec_out = 64'b1111001111010111110111110111010110111101111110111101110110011001;
          11:
            level_vec_out = 64'b1111001111010111110111110111010110111101111110111101110110011001;
          12:
            level_vec_out = 64'b1111001111010111110111110111010110111101111110111101110110111001;
          13:
            level_vec_out = 64'b1111001111010111110111110111110110111101111110111101110110111001;
          14:
            level_vec_out = 64'b1111001111010111110111110111111110111101111110111111110110111101;
          15:
            level_vec_out = 64'b1111001111010111110111110111111110111101111110111111110110111101;
          16:
            level_vec_out = 64'b1111001111010111110111110111111110111101111110111111110110111101;
          17:
            level_vec_out = 64'b1111001111010111110111110111111110111101111110111111110110111101;
          18:
            level_vec_out = 64'b1111001111010111110111110111111110111101111110111111110110111101;
          19:
            level_vec_out = 64'b1111001111010111110111110111111110111101111110111111110110111101;
          20:
            level_vec_out = 64'b1111001111010111110111111111111110111101111110111111110110111101;
          21:
            level_vec_out = 64'b1111011111010111110111111111111110111111111111111111110110111101;
          22:
            level_vec_out = 64'b1111011111010111111111111111111110111111111111111111111110111101;
          23:
            level_vec_out = 64'b1111011111010111111111111111111110111111111111111111111110111101;
          24:
            level_vec_out = 64'b1111011111010111111111111111111110111111111111111111111111111101;
          25:
            level_vec_out = 64'b1111011111010111111111111111111110111111111111111111111111111101;
          26:
            level_vec_out = 64'b1111111111010111111111111111111110111111111111111111111111111101;
          27:
            level_vec_out = 64'b1111111111010111111111111111111110111111111111111111111111111111;
          28:
            level_vec_out = 64'b1111111111010111111111111111111111111111111111111111111111111111;
          29:
            level_vec_out = 64'b1111111111010111111111111111111111111111111111111111111111111111;
          30:
            level_vec_out = 64'b1111111111011111111111111111111111111111111111111111111111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        endcase
      2:
        case (frame_id)
          0:
            level_vec_out = 64'b1011001101100100100001001011100111000111011000000011001011110101;
          1:
            level_vec_out = 64'b1011001101100100100001001011100111000111011000000011001011110101;
          2:
            level_vec_out = 64'b1011001101100100100001001011100111000111011101000011001011110101;
          3:
            level_vec_out = 64'b1011001101100100100001001011100111000111011101000011001011110101;
          4:
            level_vec_out = 64'b1011001101100100100001001011100111000111011101000011001011110101;
          5:
            level_vec_out = 64'b1011001101100100100001001011100111000111011101000011001011110101;
          6:
            level_vec_out = 64'b1011001101100100100001001011100111000111011101010011001011110101;
          7:
            level_vec_out = 64'b1011001101100100100001001011100111000111011101010011001011111101;
          8:
            level_vec_out = 64'b1011001101100100100011001011101111000111011101010011001111111101;
          9:
            level_vec_out = 64'b1011001101100100100011001011101111001111011101010011001111111101;
          10:
            level_vec_out = 64'b1011001101100100100011001011101111001111011101010011001111111101;
          11:
            level_vec_out = 64'b1011001101100100100011001011101111001111111101010011001111111101;
          12:
            level_vec_out = 64'b1011001101100100100011001011101111001111111101011011001111111101;
          13:
            level_vec_out = 64'b1011001101101100110011001011101111001111111101011011001111111101;
          14:
            level_vec_out = 64'b1011001101101100110011001011101111001111111101011011001111111101;
          15:
            level_vec_out = 64'b1011001101101100110011011011101111001111111101111011001111111101;
          16:
            level_vec_out = 64'b1111001101101100110111011011101111001111111101111011001111111101;
          17:
            level_vec_out = 64'b1111001101101110110111011011101111001111111101111011001111111101;
          18:
            level_vec_out = 64'b1111001101101110110111011011101111011111111111111011101111111101;
          19:
            level_vec_out = 64'b1111001101101110110111011011101111011111111111111011101111111101;
          20:
            level_vec_out = 64'b1111001101101110110111011011111111011111111111111011101111111101;
          21:
            level_vec_out = 64'b1111001101101110110111011011111111011111111111111011101111111101;
          22:
            level_vec_out = 64'b1111001101101110110111011011111111011111111111111011101111111101;
          23:
            level_vec_out = 64'b1111001101101111110111011011111111011111111111111011101111111101;
          24:
            level_vec_out = 64'b1111001101101111110111111011111111011111111111111011101111111101;
          25:
            level_vec_out = 64'b1111001101111111110111111011111111111111111111111011101111111101;
          26:
            level_vec_out = 64'b1111001101111111110111111011111111111111111111111011101111111101;
          27:
            level_vec_out = 64'b1111001111111111110111111011111111111111111111111011101111111111;
          28:
            level_vec_out = 64'b1111001111111111110111111111111111111111111111111011111111111111;
          29:
            level_vec_out = 64'b1111001111111111110111111111111111111111111111111011111111111111;
          30:
            level_vec_out = 64'b1111001111111111111111111111111111111111111111111011111111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111011111111111111;
        endcase
      3:
        case (frame_id)
          0:
            level_vec_out = 64'b0101000010011011010111110101010001111000111000101010101101100111;
          1:
            level_vec_out = 64'b0101000010011011010111110101010001111000111000101010101101100111;
          2:
            level_vec_out = 64'b0101000110011011010111110101010001111000111000101010101101101111;
          3:
            level_vec_out = 64'b1111000110011011010111111101010001111000111000101010101101101111;
          4:
            level_vec_out = 64'b1111000110011011010111111101010001111000111000101110101101101111;
          5:
            level_vec_out = 64'b1111000110011011010111111101110101111000111000101110101101101111;
          6:
            level_vec_out = 64'b1111000110011011010111111101110101111000111000101110101111101111;
          7:
            level_vec_out = 64'b1111000110011011010111111101110101111000111000101110101111101111;
          8:
            level_vec_out = 64'b1111001110011011010111111101111101111000111000101110101111111111;
          9:
            level_vec_out = 64'b1111001110011011011111111101111101111000111000101110101111111111;
          10:
            level_vec_out = 64'b1111011110011011111111111101111101111000111000101110101111111111;
          11:
            level_vec_out = 64'b1111011110011011111111111101111101111000111100101110101111111111;
          12:
            level_vec_out = 64'b1111011110011011111111111101111101111000111100101110101111111111;
          13:
            level_vec_out = 64'b1111011110011011111111111111111101111000111100101110101111111111;
          14:
            level_vec_out = 64'b1111011111011011111111111111111101111000111100101110101111111111;
          15:
            level_vec_out = 64'b1111011111011011111111111111111111111000111100101110101111111111;
          16:
            level_vec_out = 64'b1111011111011011111111111111111111111000111101101110101111111111;
          17:
            level_vec_out = 64'b1111011111011011111111111111111111111000111101101110101111111111;
          18:
            level_vec_out = 64'b1111011111011011111111111111111111111000111111111110101111111111;
          19:
            level_vec_out = 64'b1111011111011011111111111111111111111000111111111110101111111111;
          20:
            level_vec_out = 64'b1111011111011011111111111111111111111000111111111110101111111111;
          21:
            level_vec_out = 64'b1111011111011011111111111111111111111000111111111110101111111111;
          22:
            level_vec_out = 64'b1111011111011011111111111111111111111000111111111110101111111111;
          23:
            level_vec_out = 64'b1111011111111011111111111111111111111000111111111110101111111111;
          24:
            level_vec_out = 64'b1111111111111011111111111111111111111000111111111110101111111111;
          25:
            level_vec_out = 64'b1111111111111011111111111111111111111000111111111110101111111111;
          26:
            level_vec_out = 64'b1111111111111111111111111111111111111100111111111110101111111111;
          27:
            level_vec_out = 64'b1111111111111111111111111111111111111100111111111110101111111111;
          28:
            level_vec_out = 64'b1111111111111111111111111111111111111100111111111111111111111111;
          29:
            level_vec_out = 64'b1111111111111111111111111111111111111101111111111111111111111111;
          30:
            level_vec_out = 64'b1111111111111111111111111111111111111101111111111111111111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111101111111111111111111111111;
        endcase
      4:
        case (frame_id)
          0:
            level_vec_out = 64'b0000000101111001000100001011010001110111010001000100100110110010;
          1:
            level_vec_out = 64'b0000000101111001000100001011010001110111010001000100100110110010;
          2:
            level_vec_out = 64'b0000000101111001000100001011010001110111010001000100100110110010;
          3:
            level_vec_out = 64'b0000000101111001000100001011010001110111010001000100100110110010;
          4:
            level_vec_out = 64'b0000000101111001000100001011010001110111010001000100111110110010;
          5:
            level_vec_out = 64'b0000000101111001000100001111010001110111010001000100111110110010;
          6:
            level_vec_out = 64'b0000000101111001000100001111010001110111010001000100111110110110;
          7:
            level_vec_out = 64'b0000000101111001001100101111010001110111010001000100111110110110;
          8:
            level_vec_out = 64'b0000000101111001001100101111010001110111010001000100111110110110;
          9:
            level_vec_out = 64'b0000000101111001001100101111010001110111010001000100111111110111;
          10:
            level_vec_out = 64'b0000000101111001001100101111010001110111010001100100111111110111;
          11:
            level_vec_out = 64'b0000000101111011001100101111010001110111010001100100111111111111;
          12:
            level_vec_out = 64'b0000000101111011001100101111011001110111010001100100111111111111;
          13:
            level_vec_out = 64'b0000000101111011001100101111011001110111010001100100111111111111;
          14:
            level_vec_out = 64'b0000000101111011001100101111011011110111010001100100111111111111;
          15:
            level_vec_out = 64'b0000000101111011001100101111011011110111010001100101111111111111;
          16:
            level_vec_out = 64'b0001001101111111001100101111011011110111011001100101111111111111;
          17:
            level_vec_out = 64'b0001001101111111011100101111011011110111111001100101111111111111;
          18:
            level_vec_out = 64'b0011001101111111011100101111011011110111111001100101111111111111;
          19:
            level_vec_out = 64'b0011001111111111011100101111011011110111111011100101111111111111;
          20:
            level_vec_out = 64'b0111001111111111011100101111111011110111111011100101111111111111;
          21:
            level_vec_out = 64'b0111001111111111011100101111111011110111111011110101111111111111;
          22:
            level_vec_out = 64'b1111001111111111011101101111111011110111111011110101111111111111;
          23:
            level_vec_out = 64'b1111011111111111011101101111111111110111111011110101111111111111;
          24:
            level_vec_out = 64'b1111011111111111011101101111111111111111111011110101111111111111;
          25:
            level_vec_out = 64'b1111011111111111011101101111111111111111111011110101111111111111;
          26:
            level_vec_out = 64'b1111011111111111011101101111111111111111111011110101111111111111;
          27:
            level_vec_out = 64'b1111011111111111011101111111111111111111111011110101111111111111;
          28:
            level_vec_out = 64'b1111111111111111011101111111111111111111111011110101111111111111;
          29:
            level_vec_out = 64'b1111111111111111011101111111111111111111111111110101111111111111;
          30:
            level_vec_out = 64'b1111111111111111011101111111111111111111111111110111111111111111;
          31:
            level_vec_out = 64'b1111111111111111111101111111111111111111111111111111111111111111;
        endcase
      5:
        case (frame_id)
          0:
            level_vec_out = 64'b0100101110101000011000010010000101010011010001000110000110001000;
          1:
            level_vec_out = 64'b0100101110101000011000010010000101010011010001000110000110001000;
          2:
            level_vec_out = 64'b0100101110101000011000010010100101011011010001000110000110001000;
          3:
            level_vec_out = 64'b0100111110111000011000010010100101011011010001000110000110001000;
          4:
            level_vec_out = 64'b0100111110111000011000010010100101011011010001000110000110001000;
          5:
            level_vec_out = 64'b0100111110111000011010010010100101011011010001000110000110101000;
          6:
            level_vec_out = 64'b0100111110111000011010010010100101011011010001000110000110101000;
          7:
            level_vec_out = 64'b0100111110111000011010110010100101011111010001000110000110101000;
          8:
            level_vec_out = 64'b0100111110111000011010110010100101011111010001000110000110101000;
          9:
            level_vec_out = 64'b0100111110111001011010110010100101011111010001100110010110101000;
          10:
            level_vec_out = 64'b0110111110111001011010110011100101011111011001100110010110101000;
          11:
            level_vec_out = 64'b0110111110111001011110110011100101011111011001100110010110101000;
          12:
            level_vec_out = 64'b0110111110111001011110110011100101011111011101100111010110101000;
          13:
            level_vec_out = 64'b0110111110111001011110110011100101011111011101100111010111111000;
          14:
            level_vec_out = 64'b0110111110111001011110110011100101011111011101100111010111111000;
          15:
            level_vec_out = 64'b0110111110111001011110110011100101011111011101100111010111111000;
          16:
            level_vec_out = 64'b0110111110111001011110110011100101011111011101100111010111111000;
          17:
            level_vec_out = 64'b0110111110111001011110110011101101011111011101110111010111111001;
          18:
            level_vec_out = 64'b0111111110111001011110110011101101011111011101110111010111111001;
          19:
            level_vec_out = 64'b0111111110111011011110110011111101011111011101110111110111111001;
          20:
            level_vec_out = 64'b0111111110111011011110110011111101011111011101110111110111111001;
          21:
            level_vec_out = 64'b0111111110111011011110111011111101011111011101110111110111111001;
          22:
            level_vec_out = 64'b0111111110111111011110111011111101111111111101110111110111111001;
          23:
            level_vec_out = 64'b0111111110111111011110111011111101111111111111110111110111111001;
          24:
            level_vec_out = 64'b0111111110111111011110111011111101111111111111110111110111111001;
          25:
            level_vec_out = 64'b0111111110111111011110111011111101111111111111110111110111111011;
          26:
            level_vec_out = 64'b0111111110111111011110111011111101111111111111110111110111111011;
          27:
            level_vec_out = 64'b0111111110111111011111111011111101111111111111110111110111111011;
          28:
            level_vec_out = 64'b0111111110111111011111111011111101111111111111110111110111111111;
          29:
            level_vec_out = 64'b0111111110111111111111111011111101111111111111110111110111111111;
          30:
            level_vec_out = 64'b1111111110111111111111111011111111111111111111111111110111111111;
          31:
            level_vec_out = 64'b1111111110111111111111111011111111111111111111111111110111111111;
        endcase
      6:
        case (frame_id)
          0:
            level_vec_out = 64'b1110011111000100001001011111001001111101110011000110101001001101;
          1:
            level_vec_out = 64'b1110011111000100001011011111001001111111110011000110101001001101;
          2:
            level_vec_out = 64'b1110011111000100001011011111001001111111110011000110101001001101;
          3:
            level_vec_out = 64'b1110011111000100001011011111001011111111110011000110101001001101;
          4:
            level_vec_out = 64'b1110011111000100001011011111001011111111110011000110101001001101;
          5:
            level_vec_out = 64'b1111011111100100001011011111001011111111110011000110101001001101;
          6:
            level_vec_out = 64'b1111011111100100001011011111001011111111110011100110101001001101;
          7:
            level_vec_out = 64'b1111011111100100001011011111001011111111110011100110101001001101;
          8:
            level_vec_out = 64'b1111011111100100011111011111001011111111110011100110101001001101;
          9:
            level_vec_out = 64'b1111011111100100111111011111001011111111110011100110101001001101;
          10:
            level_vec_out = 64'b1111011111100100111111011111001011111111110011100110101001001101;
          11:
            level_vec_out = 64'b1111011111100100111111011111011011111111110011100111101001011101;
          12:
            level_vec_out = 64'b1111011111101100111111011111011011111111110011100111101101011101;
          13:
            level_vec_out = 64'b1111011111101110111111011111011011111111110011100111101101011101;
          14:
            level_vec_out = 64'b1111011111101110111111011111011011111111111011100111101101011101;
          15:
            level_vec_out = 64'b1111011111101110111111011111011011111111111011100111101111011101;
          16:
            level_vec_out = 64'b1111011111101110111111011111011011111111111011100111101111011101;
          17:
            level_vec_out = 64'b1111011111101110111111011111011011111111111011100111101111011101;
          18:
            level_vec_out = 64'b1111011111101110111111011111111011111111111011100111101111011101;
          19:
            level_vec_out = 64'b1111011111101110111111011111111011111111111011110111101111011101;
          20:
            level_vec_out = 64'b1111111111101110111111011111111111111111111011110111101111011101;
          21:
            level_vec_out = 64'b1111111111101110111111011111111111111111111011110111101111011101;
          22:
            level_vec_out = 64'b1111111111101110111111011111111111111111111011110111101111011101;
          23:
            level_vec_out = 64'b1111111111101110111111011111111111111111111011110111101111011101;
          24:
            level_vec_out = 64'b1111111111101110111111011111111111111111111011111111111111011101;
          25:
            level_vec_out = 64'b1111111111111111111111011111111111111111111011111111111111011101;
          26:
            level_vec_out = 64'b1111111111111111111111011111111111111111111011111111111111111101;
          27:
            level_vec_out = 64'b1111111111111111111111011111111111111111111011111111111111111101;
          28:
            level_vec_out = 64'b1111111111111111111111011111111111111111111011111111111111111101;
          29:
            level_vec_out = 64'b1111111111111111111111111111111111111111111011111111111111111101;
          30:
            level_vec_out = 64'b1111111111111111111111111111111111111111111011111111111111111101;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111011111111111111111101;
        endcase
      7:
        case (frame_id)
          0:
            level_vec_out = 64'b0101111110111110010111011011111110010010011011101000001111111001;
          1:
            level_vec_out = 64'b0101111110111110010111011011111110110010011011101000001111111001;
          2:
            level_vec_out = 64'b0101111110111110010111011011111110110010011011101000001111111001;
          3:
            level_vec_out = 64'b0101111110111110010111011011111110110010011011101000001111111001;
          4:
            level_vec_out = 64'b0101111110111110010111011011111110110010011111101000001111111001;
          5:
            level_vec_out = 64'b0101111110111110010111011011111110110010011111101000001111111001;
          6:
            level_vec_out = 64'b0101111110111110010111011011111110110010011111101000001111111001;
          7:
            level_vec_out = 64'b0101111110111110010111011011111110110010011111101000001111111001;
          8:
            level_vec_out = 64'b0101111110111110010111011011111110110010011111101000001111111001;
          9:
            level_vec_out = 64'b0101111110111110010111011011111110110010011111101000001111111001;
          10:
            level_vec_out = 64'b0101111110111110010111011011111110110010011111101001001111111001;
          11:
            level_vec_out = 64'b0101111110111110010111011011111110110010011111101001001111111001;
          12:
            level_vec_out = 64'b0101111110111110010111011011111110110010111111101001001111111001;
          13:
            level_vec_out = 64'b0101111110111110010111011011111110110010111111101001001111111001;
          14:
            level_vec_out = 64'b1101111110111110010111011011111110110010111111101001001111111001;
          15:
            level_vec_out = 64'b1101111110111110010111011011111110110010111111101101001111111001;
          16:
            level_vec_out = 64'b1101111110111110010111011011111110110010111111101101001111111001;
          17:
            level_vec_out = 64'b1101111110111110010111011011111110110010111111101101001111111001;
          18:
            level_vec_out = 64'b1101111110111110010111011011111110110010111111101101001111111001;
          19:
            level_vec_out = 64'b1101111110111110011111011011111110110010111111101101001111111001;
          20:
            level_vec_out = 64'b1101111110111110011111011011111110110010111111101101001111111001;
          21:
            level_vec_out = 64'b1101111110111110011111011011111110110010111111101101001111111001;
          22:
            level_vec_out = 64'b1101111110111110011111111011111110110010111111101101001111111001;
          23:
            level_vec_out = 64'b1101111110111110011111111011111110110010111111101101001111111101;
          24:
            level_vec_out = 64'b1101111110111110011111111011111110110010111111111101001111111101;
          25:
            level_vec_out = 64'b1101111110111110011111111011111110110110111111111101011111111101;
          26:
            level_vec_out = 64'b1101111110111110111111111111111110111110111111111101011111111101;
          27:
            level_vec_out = 64'b1111111110111110111111111111111110111110111111111101011111111111;
          28:
            level_vec_out = 64'b1111111110111110111111111111111110111111111111111101011111111111;
          29:
            level_vec_out = 64'b1111111111111110111111111111111111111111111111111101111111111111;
          30:
            level_vec_out = 64'b1111111111111110111111111111111111111111111111111111111111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        endcase
    endcase
  end
endmodule