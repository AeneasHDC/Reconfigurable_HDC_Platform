/**
 * @file level_hvec_gen_hdl.hpp
 * @brief This script generates HDL code for generating high-dimensional LEVEL vectors.
 * It is a novel method; for more information, please refer to our paper.
 *
 * @author Saeid Jamili and Marco Angioli
 * @note Author names are listed in alphabetical order.
 * @email <saeid.jamili@uniroma1.it>
 * @email <marco.angioli@uniroma1.it>
 *
 * @contributors
 *
 * @date Created: 24th July 2023
 * @date Last Updated: 23th August 2023
 *
 * @version 0.0.1-dev
 *
 * @institute Sapienza University of Rome
 * @cite https://doi.org/10.xxxx/yyyyy
 *
 * @section DEPENDENCIES
 * - Dependency1: Description or version details.
 * - Dependency2: Description or version details.
 *
 * @section LICENSE
 * This file is part of the Aeneas HyperCompute Platform.
 *
 * Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 *
 * @section CHANGELOG
 * @version 1.0.0-dev - 23th August 2023
 * - Initial release
 *
 * @todo
 * - Complete level vector generator function
 * - Add training
 *
 * @see
 * -
 * -
 * -
 *
 */

module level_hvec_gen #(parameter int DI_PARALLEL_W_BITS = 100) (
  input logic [3:0] frame_index,
  input logic [4:0] frame_id,
  output logic [DI_PARALLEL_W_BITS-1:0] level_vec_out
);
  always_comb begin
    case (frame_index)
      0:
        case (frame_id)
          0:
            level_vec_out = 100'b0010000100101001110010011011110101010110110101001100010001101111010101011110110011101110011000100011;
          1:
            level_vec_out = 100'b0010001100101001110010011011110101010110110101001100010001101111011101011110110011101110011000100011;
          2:
            level_vec_out = 100'b0010001100101001110010011011110101010110110101001100010001101111011101011110110011101110011000100011;
          3:
            level_vec_out = 100'b0010001100101001110010011011111101010110110101001100010001101111011101011110110011101110011000100011;
          4:
            level_vec_out = 100'b1011001100101001110110011011111101010110110101001100010001111111011101011110110011101110011000100011;
          5:
            level_vec_out = 100'b1011001100101001110110011011111101010110110101001100010001111111011101011110110011101110011000100011;
          6:
            level_vec_out = 100'b1011001100101001110110011011111101010110110101001100010001111111011101011110110011101110011000100011;
          7:
            level_vec_out = 100'b1011001100101001110110011011111101010110110101001100010001111111011101011110110011101110011000100011;
          8:
            level_vec_out = 100'b1011001100101011110110011011111101011110110101001100010001111111011101011110110011101110011000100011;
          9:
            level_vec_out = 100'b1011001100101111110110011011111101011110110101101100010101111111011101011110110011101110011000100011;
          10:
            level_vec_out = 100'b1011001100101111110110011011111101011110110101101100010101111111011111011111110111101110011000100011;
          11:
            level_vec_out = 100'b1011001100101111110110011011111101011110110101101100010101111111011111011111110111101111011000100011;
          12:
            level_vec_out = 100'b1011001100101111110110011011111101011110110101101100010111111111011111011111110111101111011010100011;
          13:
            level_vec_out = 100'b1011011100101111110110011011111101011110110101101100010111111111011111011111110111101111011010110011;
          14:
            level_vec_out = 100'b1011011100101111110110011011111101011110110101101110010111111111011111011111110111101111011011111011;
          15:
            level_vec_out = 100'b1011011110101111110110011011111111011110110101101110010111111111011111011111110111101111011011111011;
          16:
            level_vec_out = 100'b1011011110101111110110011011111111011110110101101110010111111111011111011111111111111111011011111011;
          17:
            level_vec_out = 100'b1011011110101111110110011011111111011110110101101110010111111111011111011111111111111111011011111011;
          18:
            level_vec_out = 100'b1011011110111111110110011011111111011110110101101110010111111111011111011111111111111111011011111011;
          19:
            level_vec_out = 100'b1011011110111111110110011011111111011110110101101110010111111111011111011111111111111111011011111111;
          20:
            level_vec_out = 100'b1011011110111111110110111111111111011110110101101110010111111111011111011111111111111111011011111111;
          21:
            level_vec_out = 100'b1011011110111111110110111111111111011110110101111110010111111111111111011111111111111111011011111111;
          22:
            level_vec_out = 100'b1011011110111111111110111111111111011110110101111110010111111111111111111111111111111111011011111111;
          23:
            level_vec_out = 100'b1011011111111111111110111111111111011110110101111110010111111111111111111111111111111111011011111111;
          24:
            level_vec_out = 100'b1011011111111111111111111111111111011110110111111110010111111111111111111111111111111111011011111111;
          25:
            level_vec_out = 100'b1011011111111111111111111111111111011110110111111110011111111111111111111111111111111111011011111111;
          26:
            level_vec_out = 100'b1011111111111111111111111111111111011111110111111110011111111111111111111111111111111111011011111111;
          27:
            level_vec_out = 100'b1011111111111111111111111111111111011111110111111110011111111111111111111111111111111111111111111111;
          28:
            level_vec_out = 100'b1111111111111111111111111111111111011111110111111110011111111111111111111111111111111111111111111111;
          29:
            level_vec_out = 100'b1111111111111111111111111111111111011111110111111110011111111111111111111111111111111111111111111111;
        endcase
      1:
        case (frame_id)
          0:
            level_vec_out = 100'b1010001101100110111000001000010110011000111010010010110010100100111011000010011111001001000100111111;
          1:
            level_vec_out = 100'b1010001111100110111000001000010110011000111010010110110010100100111011000010011111001001000100111111;
          2:
            level_vec_out = 100'b1010101111100110111000001000010110011000111010010110110110100100111111000010011111001001000100111111;
          3:
            level_vec_out = 100'b1010101111100110111000001000010110011000111110010110110110100100111111000010011111001001001100111111;
          4:
            level_vec_out = 100'b1010101111100110111000001000010110011000111110010110110110100100111111000010011111001001001100111111;
          5:
            level_vec_out = 100'b1010101111100110111100001000110110011000111110010110110110100100111111000010011111001001001100111111;
          6:
            level_vec_out = 100'b1010101111100110111100001010111110011000111110010110110110100100111111000011011111001001001100111111;
          7:
            level_vec_out = 100'b1010101111100110111100101010111110011000111110010110110110100100111111000011011111001001001100111111;
          8:
            level_vec_out = 100'b1010101111100110111100101010111110011000111110010110110110100100111111000011011111001001001100111111;
          9:
            level_vec_out = 100'b1010101111100110111100101010111110011000111110010110110110100100111111010011011111001011001100111111;
          10:
            level_vec_out = 100'b1010101111100110111100101010111110011000111110010110110110100100111111010011011111001011001110111111;
          11:
            level_vec_out = 100'b1010101111100110111100101010111110011000111110010110110110100100111111010011011111001011001110111111;
          12:
            level_vec_out = 100'b1110101111100110111100101010111110011000111110010110110110100100111111010111011111001011001110111111;
          13:
            level_vec_out = 100'b1110101111100110111100101011111110011000111111010110110110100100111111010111011111001111001110111111;
          14:
            level_vec_out = 100'b1110101111100110111100101011111110011000111111010110110110100100111111010111111111001111001110111111;
          15:
            level_vec_out = 100'b1110101111100110111100101011111110011000111111010110110110101100111111010111111111101111001110111111;
          16:
            level_vec_out = 100'b1110101111100110111100101011111110011001111111010110110110101100111111010111111111101111001110111111;
          17:
            level_vec_out = 100'b1110101111100110111101101011111110011011111111010110110110101100111111010111111111101111001110111111;
          18:
            level_vec_out = 100'b1110111111100110111101101011111110011011111111010110111110101100111111010111111111101111101110111111;
          19:
            level_vec_out = 100'b1110111111100111111101101011111110011011111111010110111110101100111111010111111111111111101110111111;
          20:
            level_vec_out = 100'b1110111111111111111101101011111110011011111111010110111110101100111111010111111111111111111110111111;
          21:
            level_vec_out = 100'b1111111111111111111101111011111111011011111111110110111110101100111111010111111111111111111110111111;
          22:
            level_vec_out = 100'b1111111111111111111101111011111111011011111111110110111110101100111111010111111111111111111110111111;
          23:
            level_vec_out = 100'b1111111111111111111101111111111111011011111111110110111110111100111111010111111111111111111110111111;
          24:
            level_vec_out = 100'b1111111111111111111101111111111111011011111111110110111110111100111111010111111111111111111110111111;
          25:
            level_vec_out = 100'b1111111111111111111101111111111111011011111111110111111110111111111111010111111111111111111110111111;
          26:
            level_vec_out = 100'b1111111111111111111111111111111111111011111111110111111110111111111111110111111111111111111111111111;
          27:
            level_vec_out = 100'b1111111111111111111111111111111111111011111111110111111111111111111111110111111111111111111111111111;
          28:
            level_vec_out = 100'b1111111111111111111111111111111111111011111111110111111111111111111111110111111111111111111111111111;
          29:
            level_vec_out = 100'b1111111111111111111111111111111111111011111111110111111111111111111111110111111111111111111111111111;
        endcase
      2:
        case (frame_id)
          0:
            level_vec_out = 100'b0001001101001000100111001111111000000100110111110111101011110010100000001001100001111111011101110100;
          1:
            level_vec_out = 100'b0001101101001000100111001111111000000100111111110111101011110010100000001001100001111111011101110100;
          2:
            level_vec_out = 100'b0001101101001000100111001111111000000100111111110111101011110010100000001001100001111111011101110100;
          3:
            level_vec_out = 100'b0001101101001000100111001111111000000100111111110111101011110010100000001001100001111111011101110100;
          4:
            level_vec_out = 100'b0001101101001000110111001111111000000100111111110111101011110010100000001001100001111111011101110100;
          5:
            level_vec_out = 100'b0001111101001000110111001111111010000100111111110111101011110010100000001001100001111111011101110100;
          6:
            level_vec_out = 100'b0001111101001000110111001111111010000100111111110111101011110010100000001001100001111111011101110100;
          7:
            level_vec_out = 100'b0001111111001000110111001111111011100100111111110111101011110010100000001001100001111111011101110100;
          8:
            level_vec_out = 100'b0011111111001000110111001111111011100101111111110111101011110010100000001001100001111111011101110100;
          9:
            level_vec_out = 100'b0011111111001010110111001111111011100101111111110111101011110010100000001101100001111111011101110100;
          10:
            level_vec_out = 100'b0011111111001010111111001111111011100101111111110111101011110010100000001101100001111111011101110100;
          11:
            level_vec_out = 100'b1011111111001010111111001111111011100101111111110111101011110010100001001101100001111111011101110100;
          12:
            level_vec_out = 100'b1011111111001010111111001111111011100101111111111111101011110010100001001101100001111111011101110110;
          13:
            level_vec_out = 100'b1011111111001010111111001111111111100101111111111111101011110010100001001101100001111111011101110110;
          14:
            level_vec_out = 100'b1011111111001010111111001111111111100111111111111111101011110010100011001111100001111111011101110110;
          15:
            level_vec_out = 100'b1011111111001010111111001111111111110111111111111111101011110110100011101111100001111111011101111110;
          16:
            level_vec_out = 100'b1011111111011010111111001111111111110111111111111111101011110110100011101111100001111111011101111110;
          17:
            level_vec_out = 100'b1011111111011010111111001111111111110111111111111111101011110110100011101111100001111111011101111110;
          18:
            level_vec_out = 100'b1011111111011010111111101111111111110111111111111111101011110110100011101111100001111111011101111110;
          19:
            level_vec_out = 100'b1011111111011010111111101111111111110111111111111111101011110110100011101111100001111111011101111110;
          20:
            level_vec_out = 100'b1011111111011010111111101111111111111111111111111111101011110110110011101111100011111111011101111110;
          21:
            level_vec_out = 100'b1011111111011010111111101111111111111111111111111111101011110110110011111111100011111111011101111110;
          22:
            level_vec_out = 100'b1111111111111010111111101111111111111111111111111111101011110110110011111111101011111111011101111110;
          23:
            level_vec_out = 100'b1111111111111010111111101111111111111111111111111111101011110110110011111111101011111111011101111110;
          24:
            level_vec_out = 100'b1111111111111110111111101111111111111111111111111111111011110110110011111111101011111111011101111110;
          25:
            level_vec_out = 100'b1111111111111111111111101111111111111111111111111111111011110110111011111111101011111111011111111111;
          26:
            level_vec_out = 100'b1111111111111111111111101111111111111111111111111111111011111110111011111111101011111111011111111111;
          27:
            level_vec_out = 100'b1111111111111111111111101111111111111111111111111111111011111110111011111111101011111111011111111111;
          28:
            level_vec_out = 100'b1111111111111111111111101111111111111111111111111111111011111110111011111111111011111111011111111111;
          29:
            level_vec_out = 100'b1111111111111111111111101111111111111111111111111111111011111111111011111111111011111111111111111111;
        endcase
      3:
        case (frame_id)
          0:
            level_vec_out = 100'b1111110011001010010011100111111011000101101000010000100101010111011101101011110101001001011000010101;
          1:
            level_vec_out = 100'b1111110011011010010011100111111011000101101000010010100101010111011101101011110101001001011000010101;
          2:
            level_vec_out = 100'b1111110011011010010011100111111011000101101000010010100101010111011101111011110111001001011000010101;
          3:
            level_vec_out = 100'b1111110011011010010011100111111011000101101000010010100101010111011101111011110111001001011000010101;
          4:
            level_vec_out = 100'b1111110011011010010011100111111011000101101000010010100101010111011101111011110111001111011000010101;
          5:
            level_vec_out = 100'b1111110011011010010011100111111011000101101000010010100101010111011101111011110111001111011000010101;
          6:
            level_vec_out = 100'b1111110011011010010011101111111011000101111000010010100101010111011101111011110111001111011000010101;
          7:
            level_vec_out = 100'b1111110011011010010011101111111011000101111000010010100101010111011101111011110111001111011000010101;
          8:
            level_vec_out = 100'b1111110011011010010011111111111011000101111000010010100101010111011101111011110111011111011000010101;
          9:
            level_vec_out = 100'b1111110011011010010011111111111011000101111000010010100101011111011101111011110111011111011000010101;
          10:
            level_vec_out = 100'b1111110111011010010011111111111011000101111000010010100101011111011101111011110111011111011000010101;
          11:
            level_vec_out = 100'b1111110111011010010011111111111011001111111000010010100101011111011101111011110111011111011000010101;
          12:
            level_vec_out = 100'b1111111111011010010011111111111011001111111000010010100101011111011111111011110111011111011000010101;
          13:
            level_vec_out = 100'b1111111111011010010011111111111011001111111000011010100101011111011111111011110111011111011000010101;
          14:
            level_vec_out = 100'b1111111111011010010011111111111011001111111000011010100101011111011111111011111111011111011000010111;
          15:
            level_vec_out = 100'b1111111111011010010011111111111011001111111000011010100101011111011111111011111111011111011000010111;
          16:
            level_vec_out = 100'b1111111111011010010011111111111011001111111000011010100101011111011111111011111111011111011000110111;
          17:
            level_vec_out = 100'b1111111111011010110011111111111011001111111000011011110101011111011111111011111111011111011000110111;
          18:
            level_vec_out = 100'b1111111111011110110011111111111011001111111000011011110101011111011111111011111111011111111000110111;
          19:
            level_vec_out = 100'b1111111111011110111111111111111011001111111000011011110101011111011111111011111111011111111000111111;
          20:
            level_vec_out = 100'b1111111111011110111111111111111111001111111000011011110111111111011111111011111111011111111010111111;
          21:
            level_vec_out = 100'b1111111111011111111111111111111111001111111000011011110111111111111111111011111111011111111010111111;
          22:
            level_vec_out = 100'b1111111111011111111111111111111111001111111000011011110111111111111111111011111111011111111010111111;
          23:
            level_vec_out = 100'b1111111111111111111111111111111111001111111000011011110111111111111111111011111111011111111010111111;
          24:
            level_vec_out = 100'b1111111111111111111111111111111111001111111001011011110111111111111111111011111111011111111010111111;
          25:
            level_vec_out = 100'b1111111111111111111111111111111111101111111001011011110111111111111111111011111111011111111010111111;
          26:
            level_vec_out = 100'b1111111111111111111111111111111111101111111001011011110111111111111111111011111111011111111010111111;
          27:
            level_vec_out = 100'b1111111111111111111111111111111111111111111011011011110111111111111111111011111111011111111010111111;
          28:
            level_vec_out = 100'b1111111111111111111111111111111111111111111011111111110111111111111111111011111111111111111010111111;
          29:
            level_vec_out = 100'b1111111111111111111111111111111111111111111011111111110111111111111111111111111111111111111011111111;
        endcase
      4:
        case (frame_id)
          0:
            level_vec_out = 100'b0001111110100001010100000110110101000001010111001000000011011010101111100001110101001111110000101100;
          1:
            level_vec_out = 100'b0001111110100001010100000110110101000001010111001000000011011010101111100001110111001111110000101100;
          2:
            level_vec_out = 100'b0001111110100001010100000110110101100001010111001000000011011010101111100001110111001111110000101110;
          3:
            level_vec_out = 100'b0001111110100001010100000110110101100001110111001000000111011010101111100001110111001111110010101110;
          4:
            level_vec_out = 100'b0001111110100001010100100111110101100001110111001000000111011010101111100001110111001111110010101110;
          5:
            level_vec_out = 100'b0001111110110001010100100111110101100001110111001000000111011010101111100001110111001111110010101110;
          6:
            level_vec_out = 100'b0001111110110001010100100111110101100001110111001000100111011011101111100001110111001111110010101110;
          7:
            level_vec_out = 100'b0001111110110001010100100111110101100001110111001000100111011011101111110001110111001111110010101110;
          8:
            level_vec_out = 100'b0001111110110001010100100111110101100011110111001000100111011011101111111001110111001111110010101110;
          9:
            level_vec_out = 100'b0001111110110001010100100111110101100011110111001000100111011011111111111001110111001111111010101110;
          10:
            level_vec_out = 100'b0001111110110001010100100111110101100011110111001000100111011011111111111001110111001111111010101110;
          11:
            level_vec_out = 100'b0001111110110001010100100111110101100011110111001000100111011011111111111001110111001111111010101110;
          12:
            level_vec_out = 100'b0001111110110001010100100111110101100011110111001000100111011011111111111001110111001111111010101110;
          13:
            level_vec_out = 100'b0001111110110001010100100111110101100011110111001010100111011011111111111001110111001111111010101110;
          14:
            level_vec_out = 100'b0001111110111001010100100111110101100011110111001010100111011011111111111001110111001111111010101110;
          15:
            level_vec_out = 100'b0001111110111001010100100111110101100011110111001010100111011011111111111001110111001111111010101110;
          16:
            level_vec_out = 100'b0001111110111001110110100111110101100011110111101010100111011011111111111001110111001111111010101110;
          17:
            level_vec_out = 100'b0001111110111001110110100111110101100011110111101010100111011011111111111001110111001111111011101110;
          18:
            level_vec_out = 100'b0001111111111001111110100111110101100011110111101010100111011011111111111001110111001111111011101110;
          19:
            level_vec_out = 100'b0001111111111001111110101111110101100011110111101010100111011011111111111001110111001111111011101110;
          20:
            level_vec_out = 100'b0001111111111001111110101111110101110011110111101010100111011011111111111001110111001111111011101110;
          21:
            level_vec_out = 100'b0101111111111001111110111111110111110011110111101110100111011011111111111001110111001111111011101110;
          22:
            level_vec_out = 100'b0101111111111001111110111111111111110011111111101110100111011011111111111101110111001111111011101110;
          23:
            level_vec_out = 100'b0101111111111001111111111111111111110011111111101110100111011011111111111101110111001111111011101111;
          24:
            level_vec_out = 100'b0101111111111001111111111111111111111011111111101111100111011111111111111101110111001111111011111111;
          25:
            level_vec_out = 100'b0101111111111001111111111111111111111011111111101111100111011111111111111101110111001111111011111111;
          26:
            level_vec_out = 100'b0101111111111101111111111111111111111011111111101111100111011111111111111101110111011111111011111111;
          27:
            level_vec_out = 100'b0101111111111111111111111111111111111011111111101111100111011111111111111101110111011111111011111111;
          28:
            level_vec_out = 100'b1111111111111111111111111111111111111011111111101111101111011111111111111101110111011111111011111111;
          29:
            level_vec_out = 100'b1111111111111111111111111111111111111111111111101111101111011111111111111101111111011111111011111111;
        endcase
      5:
        case (frame_id)
          0:
            level_vec_out = 100'b0111011001010010000011111000000000111001011000001111100110100100010011100101101110000100111110110111;
          1:
            level_vec_out = 100'b0111011001010010000011111100000000111001011000001111100110100100010011100101101110000100111110110111;
          2:
            level_vec_out = 100'b0111011001010010000011111100000000111001011000001111100110100100110011100101101110000100111110110111;
          3:
            level_vec_out = 100'b0111011001010010000011111100000000111001011100101111100110100100110011100101101110000100111110110111;
          4:
            level_vec_out = 100'b0111011001010010000011111100001000111001011110101111100110100100110011100101101110000100111110110111;
          5:
            level_vec_out = 100'b0111011001110010000011111100001000111001011110101111100110100100110011100101101110000100111110110111;
          6:
            level_vec_out = 100'b0111011001110010000011111100001000111001011110101111100110110100110011110101101110000100111110110111;
          7:
            level_vec_out = 100'b0111011001110010000011111100001000111001011110101111100110110100110011110101101110000100111110110111;
          8:
            level_vec_out = 100'b0111011001110010000011111100001000111011011110101111100110110100110011110101101110100100111110110111;
          9:
            level_vec_out = 100'b0111011001110110000011111100001000111011011111101111100110110100110011110101101110100100111110110111;
          10:
            level_vec_out = 100'b0111011001110110000011111100101000111011011111101111100111110100110011110111101110100100111110110111;
          11:
            level_vec_out = 100'b0111011001111110100011111100101000111011011111101111100111110100110011110111101110100100111110110111;
          12:
            level_vec_out = 100'b0111011001111110100011111100101001111011011111101111100111110100110011110111101110100110111110111111;
          13:
            level_vec_out = 100'b0111011001111110110011111100101001111011011111101111100111111100110011110111101110100110111110111111;
          14:
            level_vec_out = 100'b0111011001111110110011111100101001111011011111101111100111111100110011110111101110100110111111111111;
          15:
            level_vec_out = 100'b0111011001111110110011111101101001111011011111101111110111111100110011110111101110100110111111111111;
          16:
            level_vec_out = 100'b0111011001111110110011111101101001111011011111111111110111111100110011110111111110100110111111111111;
          17:
            level_vec_out = 100'b0111011001111110110011111101101001111011011111111111110111111101110011110111111110100110111111111111;
          18:
            level_vec_out = 100'b0111011001111110110011111101101001111011011111111111110111111101110011111111111110101110111111111111;
          19:
            level_vec_out = 100'b0111011001111110110011111111101001111011111111111111110111111101111011111111111110101110111111111111;
          20:
            level_vec_out = 100'b0111011001111110110011111111101001111011111111111111110111111101111011111111111110101110111111111111;
          21:
            level_vec_out = 100'b0111011001111110110011111111101001111011111111111111110111111101111011111111111110101110111111111111;
          22:
            level_vec_out = 100'b0111011001111110110011111111101111111011111111111111110111111101111011111111111110101110111111111111;
          23:
            level_vec_out = 100'b0111011001111110110011111111101111111011111111111111110111111101111011111111111110101110111111111111;
          24:
            level_vec_out = 100'b0111011001111110110011111111101111111011111111111111110111111101111011111111111110101110111111111111;
          25:
            level_vec_out = 100'b0111011101111110111011111111101111111011111111111111110111111101111011111111111110101110111111111111;
          26:
            level_vec_out = 100'b1111011101111110111011111111101111111011111111111111110111111101111011111111111110101111111111111111;
          27:
            level_vec_out = 100'b1111011101111111111111111111111111111011111111111111110111111101111011111111111110101111111111111111;
          28:
            level_vec_out = 100'b1111011111111111111111111111111111111011111111111111110111111101111011111111111110101111111111111111;
          29:
            level_vec_out = 100'b1111011111111111111111111111111111111011111111111111111111111101111011111111111110111111111111111111;
        endcase
      6:
        case (frame_id)
          0:
            level_vec_out = 100'b0000000101011011110010100011111010110001010101000101100001001011001001011000111110001110111001110000;
          1:
            level_vec_out = 100'b0000000101011011110010100111111010110001010101100101100001101011001001011000111110001110111001110000;
          2:
            level_vec_out = 100'b0000000101011011110010100111111010110001010101100101100001101011001001011000111110001110111001110100;
          3:
            level_vec_out = 100'b0000000101011011110010100111111010110001010101100101100001101011001001011000111110101111111001110100;
          4:
            level_vec_out = 100'b0000000101011011110110100111111010110001010101100101100001101011001001011000111110101111111011110100;
          5:
            level_vec_out = 100'b1000000101011011110110100111111010110001010101100101100001101011001001011000111110101111111011110100;
          6:
            level_vec_out = 100'b1000000101011111110110100111111010110001010101100101100001101011001001011000111110101111111011110110;
          7:
            level_vec_out = 100'b1010000101011111110110100111111010110001010101100101101001111011101001011000111110101111111011110110;
          8:
            level_vec_out = 100'b1010000101011111110110100111111010110001010101100101101001111011101001011000111110101111111011110110;
          9:
            level_vec_out = 100'b1010000101011111110110100111111010110001010101110101111001111011101001011000111110101111111011110110;
          10:
            level_vec_out = 100'b1010000101011111110110100111111010110001010101110101111001111011101001011000111110101111111011110110;
          11:
            level_vec_out = 100'b1010000101011111110110100111111110110001010101110101111001111011101001011010111110101111111011110110;
          12:
            level_vec_out = 100'b1011000101011111110110100111111110110001010101110101111001111011101001011010111110101111111111110110;
          13:
            level_vec_out = 100'b1011000101011111110111100111111110110001010111110101111001111011101001011010111110101111111111111110;
          14:
            level_vec_out = 100'b1011000101011111110111100111111110110001010111110101111001111011101001011010111110111111111111111110;
          15:
            level_vec_out = 100'b1011000101011111110111100111111110110001010111110101111001111011111001011010111110111111111111111110;
          16:
            level_vec_out = 100'b1011000101011111110111100111111110110001010111110101111011111011111001011010111110111111111111111110;
          17:
            level_vec_out = 100'b1011000101011111110111100111111110111001011111110101111011111011111001011010111110111111111111111110;
          18:
            level_vec_out = 100'b1011000101011111110111100111111110111001011111110101111011111011111001011010111110111111111111111110;
          19:
            level_vec_out = 100'b1011100101011111110111100111111110111001011111111101111011111011111011011010111111111111111111111110;
          20:
            level_vec_out = 100'b1011100101011111110111100111111110111101011111111101111011111011111011011010111111111111111111111110;
          21:
            level_vec_out = 100'b1011100101011111110111100111111110111101111111111101111011111011111011011010111111111111111111111110;
          22:
            level_vec_out = 100'b1011100101011111110111100111111111111101111111111101111011111011111011011010111111111111111111111110;
          23:
            level_vec_out = 100'b1011100101011111110111111111111111111101111111111101111011111011111111011010111111111111111111111110;
          24:
            level_vec_out = 100'b1011110101111111111111111111111111111101111111111101111011111011111111011011111111111111111111111110;
          25:
            level_vec_out = 100'b1011111101111111111111111111111111111101111111111101111011111011111111011011111111111111111111111110;
          26:
            level_vec_out = 100'b1111111101111111111111111111111111111101111111111101111011111011111111011011111111111111111111111110;
          27:
            level_vec_out = 100'b1111111111111111111111111111111111111101111111111111111011111011111111011011111111111111111111111110;
          28:
            level_vec_out = 100'b1111111111111111111111111111111111111101111111111111111011111111111111011011111111111111111111111110;
          29:
            level_vec_out = 100'b1111111111111111111111111111111111111101111111111111111011111111111111111111111111111111111111111111;
        endcase
      7:
        case (frame_id)
          0:
            level_vec_out = 100'b1001001110011010111111001011011111010001100011011100101011110110011000111010010011000010000111011100;
          1:
            level_vec_out = 100'b1001001110011010111111001011011111010001101011011100101011110110011000111010010011000010000111011100;
          2:
            level_vec_out = 100'b1001101110011010111111001011011111010001101011011100101011110110011000111010010011000011001111011100;
          3:
            level_vec_out = 100'b1001101110011010111111001011011111011001101011011100101011110110011000111010010011000011001111011100;
          4:
            level_vec_out = 100'b1001101110011010111111001011011111011001101011011100101011110110111000111010010011000011001111011100;
          5:
            level_vec_out = 100'b1101101110011010111111001011011111011011101011011100101011110110111000111010010011000011001111011100;
          6:
            level_vec_out = 100'b1101101110011010111111001011011111011011101011011100101011110110111000111110010011000011001111011101;
          7:
            level_vec_out = 100'b1101101110011010111111001011011111011011101011011100101011110110111000111110010011000011001111011101;
          8:
            level_vec_out = 100'b1101101110011010111111001011011111011011101011011100101011110110111000111110110011010011001111011101;
          9:
            level_vec_out = 100'b1101101110011010111111001011011111011011101011011100101011110110111000111110110011010011001111011101;
          10:
            level_vec_out = 100'b1101101110011010111111001011011111011011101011011100101011110110111000111110110011010111001111011101;
          11:
            level_vec_out = 100'b1111101110011010111111001011011111011011101011011100111011110110111000111110110011010111001111011101;
          12:
            level_vec_out = 100'b1111101110011010111111001011011111011011101011011100111011110110111000111110110011010111001111011101;
          13:
            level_vec_out = 100'b1111101110011010111111001011011111011011101011011100111011110110111000111110110011010111001111011101;
          14:
            level_vec_out = 100'b1111101110011010111111001011011111011011101011011100111011110110111000111111110011010111001111011101;
          15:
            level_vec_out = 100'b1111101110011011111111001011111111011011101011011100111011111110111000111111111011010111001111011101;
          16:
            level_vec_out = 100'b1111101111011011111111001011111111011011101011111100111011111110111000111111111011010111001111011101;
          17:
            level_vec_out = 100'b1111101111011011111111001011111111111011101011111100111011111110111000111111111011010111011111011101;
          18:
            level_vec_out = 100'b1111101111011011111111001011111111111011101011111100111011111110111001111111111011110111011111011101;
          19:
            level_vec_out = 100'b1111101111011011111111001011111111111011101011111100111011111110111001111111111011110111011111011101;
          20:
            level_vec_out = 100'b1111101111011011111111001011111111111011101011111100111011111110111001111111111011110111011111011101;
          21:
            level_vec_out = 100'b1111101111011011111111001011111111111011101011111100111011111110111001111111111011110111011111011101;
          22:
            level_vec_out = 100'b1111101111011011111111001111111111111011101011111111111011111110111001111111111011110111011111011101;
          23:
            level_vec_out = 100'b1111101111011011111111001111111111111011101011111111111011111110111101111111111011110111011111011111;
          24:
            level_vec_out = 100'b1111101111011011111111001111111111111011101011111111111011111110111101111111111011110111011111011111;
          25:
            level_vec_out = 100'b1111111111011011111111001111111111111111101011111111111111111110111101111111111011110111011111011111;
          26:
            level_vec_out = 100'b1111111111011011111111101111111111111111101011111111111111111110111111111111111011110111011111011111;
          27:
            level_vec_out = 100'b1111111111011011111111101111111111111111101011111111111111111110111111111111111111110111111111111111;
          28:
            level_vec_out = 100'b1111111111011111111111111111111111111111111011111111111111111110111111111111111111111111111111111111;
          29:
            level_vec_out = 100'b1111111111011111111111111111111111111111111111111111111111111110111111111111111111111111111111111111;
        endcase
      8:
        case (frame_id)
          0:
            level_vec_out = 100'b1011111100101010110101100010000001001000011001000110101101011101111001010100110101010100111100100000;
          1:
            level_vec_out = 100'b1011111100101010110101100010001101001000011001000110101101011101111001010100110101010100111100100000;
          2:
            level_vec_out = 100'b1011111100101011110101100010001101001000011001000110101101011101111001010100110101010100111100100100;
          3:
            level_vec_out = 100'b1111111100101011110101100010001101001000011001010110101101011101111001010100110101010101111110100100;
          4:
            level_vec_out = 100'b1111111100101011110101100010001101001000011001010110101101011101111001010100110101010101111110100100;
          5:
            level_vec_out = 100'b1111111100101011110101100010001101001000011001110110101101011101111011010100110101011101111110100101;
          6:
            level_vec_out = 100'b1111111100101011110101100010001101101000111001110110101101011101111011010101110101011101111110100101;
          7:
            level_vec_out = 100'b1111111100101011110101110010001101101010111001110110101101011101111011010101111101011101111110100101;
          8:
            level_vec_out = 100'b1111111100101011110101110010001101101010111001110110101101011101111011010101111101011101111110100101;
          9:
            level_vec_out = 100'b1111111100101011110101110010001111101010111001110110101101011101111111010101111101011101111110100101;
          10:
            level_vec_out = 100'b1111111100101011111101110010001111101010111001110110101101011101111111010101111101111101111110100101;
          11:
            level_vec_out = 100'b1111111100101011111101110010001111101010111011110110101101011101111111010101111101111111111110110101;
          12:
            level_vec_out = 100'b1111111100101011111111110010001111101010111011110111101101011101111111010101111101111111111110110101;
          13:
            level_vec_out = 100'b1111111100101011111111110010001111101010111011110111101101011111111111010101111101111111111110110101;
          14:
            level_vec_out = 100'b1111111100101011111111110010001111101010111111111111101101011111111111010101111101111111111110111101;
          15:
            level_vec_out = 100'b1111111100101011111111110010001111101010111111111111101101011111111111010101111101111111111110111101;
          16:
            level_vec_out = 100'b1111111100101011111111110010001111101010111111111111101101011111111111010101111101111111111110111101;
          17:
            level_vec_out = 100'b1111111100101011111111110010001111101010111111111111101101011111111111010101111101111111111110111101;
          18:
            level_vec_out = 100'b1111111100101011111111110010001111101010111111111111101101011111111111010111111101111111111110111111;
          19:
            level_vec_out = 100'b1111111100101011111111110010001111101010111111111111101101111111111111010111111101111111111110111111;
          20:
            level_vec_out = 100'b1111111110101011111111110010001111101010111111111111101101111111111111010111111101111111111110111111;
          21:
            level_vec_out = 100'b1111111110101011111111110010001111101010111111111111101101111111111111010111111111111111111110111111;
          22:
            level_vec_out = 100'b1111111111101011111111110110001111101010111111111111101101111111111111010111111111111111111110111111;
          23:
            level_vec_out = 100'b1111111111101011111111110110101111101010111111111111101101111111111111011111111111111111111110111111;
          24:
            level_vec_out = 100'b1111111111111011111111110110101111101010111111111111101101111111111111011111111111111111111111111111;
          25:
            level_vec_out = 100'b1111111111111011111111110110101111101011111111111111101101111111111111011111111111111111111111111111;
          26:
            level_vec_out = 100'b1111111111111011111111110110101111101011111111111111101101111111111111011111111111111111111111111111;
          27:
            level_vec_out = 100'b1111111111111111111111110111101111101011111111111111101101111111111111011111111111111111111111111111;
          28:
            level_vec_out = 100'b1111111111111111111111110111111111101011111111111111101101111111111111011111111111111111111111111111;
          29:
            level_vec_out = 100'b1111111111111111111111111111111111111011111111111111111101111111111111011111111111111111111111111111;
        endcase
      9:
        case (frame_id)
          0:
            level_vec_out = 100'b1110100011101100000111011100000100110101100000010101010010010110101110011111101110010010010110001101;
          1:
            level_vec_out = 100'b1110100011101100000111011100000100110101100000010101010010010110101110011111101110010010010110001101;
          2:
            level_vec_out = 100'b1110100011111100000111011100000100111101100000010101010010010110101110011111101110010010010110001101;
          3:
            level_vec_out = 100'b1110100011111100000111011100000110111101100000010101010010010110101110011111101110010010010110001101;
          4:
            level_vec_out = 100'b1110100011111100000111011100000110111111100000010101010010010110101110011111101111010010010110001101;
          5:
            level_vec_out = 100'b1110100011111100000111111100000110111111100000010111010010010110101110011111101111010010010110011101;
          6:
            level_vec_out = 100'b1110100011111100000111111100000110111111100000010111010010010110101110011111101111010010010110011101;
          7:
            level_vec_out = 100'b1110100011111100100111111101000110111111100100010111010010010110101111011111101111010010010110011101;
          8:
            level_vec_out = 100'b1110100011111100100111111101001110111111100110010111011010010110101111011111111111010010010110011101;
          9:
            level_vec_out = 100'b1110100011111100100111111101001110111111100110010111011010010110101111011111111111010010010110011101;
          10:
            level_vec_out = 100'b1110101011111110100111111101001111111111100110010111011010010110101111011111111111010010110110011101;
          11:
            level_vec_out = 100'b1110101011111111100111111101101111111111100110010111011010010110101111011111111111010010110110011101;
          12:
            level_vec_out = 100'b1110101011111111100111111111101111111111100110010111011010010110101111011111111111010010110110011101;
          13:
            level_vec_out = 100'b1110101111111111110111111111101111111111100110010111011010010110101111011111111111010010110110011101;
          14:
            level_vec_out = 100'b1110101111111111110111111111101111111111100110010111011010010110101111011111111111010010110110011101;
          15:
            level_vec_out = 100'b1110101111111111110111111111101111111111100110010111011010010110101111011111111111010110110110011101;
          16:
            level_vec_out = 100'b1110111111111111110111111111101111111111110110010111011010010110101111011111111111010111110110011101;
          17:
            level_vec_out = 100'b1111111111111111110111111111101111111111110110010111011010010110101111011111111111011111111111111101;
          18:
            level_vec_out = 100'b1111111111111111110111111111101111111111110110010111011010010110111111011111111111011111111111111101;
          19:
            level_vec_out = 100'b1111111111111111110111111111101111111111110110010111011010010110111111011111111111111111111111111101;
          20:
            level_vec_out = 100'b1111111111111111110111111111101111111111110110010111111010010110111111011111111111111111111111111101;
          21:
            level_vec_out = 100'b1111111111111111110111111111101111111111110110010111111010110110111111011111111111111111111111111101;
          22:
            level_vec_out = 100'b1111111111111111110111111111101111111111110110010111111010110110111111011111111111111111111111111101;
          23:
            level_vec_out = 100'b1111111111111111110111111111101111111111110110010111111111110111111111011111111111111111111111111101;
          24:
            level_vec_out = 100'b1111111111111111110111111111101111111111110111010111111111110111111111011111111111111111111111111101;
          25:
            level_vec_out = 100'b1111111111111111110111111111101111111111110111010111111111110111111111011111111111111111111111111101;
          26:
            level_vec_out = 100'b1111111111111111111111111111101111111111110111010111111111111111111111011111111111111111111111111101;
          27:
            level_vec_out = 100'b1111111111111111111111111111101111111111110111010111111111111111111111011111111111111111111111111101;
          28:
            level_vec_out = 100'b1111111111111111111111111111111111111111110111010111111111111111111111011111111111111111111111111101;
          29:
            level_vec_out = 100'b1111111111111111111111111111111111111111110111010111111111111111111111111111111111111111111111111101;
        endcase
    endcase
  end
endmodule