
/**
 * @file class_hvec_gen_hdl.hpp
 * @brief This script generates HDL code for generating high-dimensional class vectors.
 * It is a novel method; for more information, please refer to our paper.
 *
 * @author Saeid Jamili and Marco Angioli
 * @note Author names are listed in alphabetical order.
 * @email <saeid.jamili@uniroma1.it>
 * @email <marco.angioli@uniroma1.it>
 *
 * @contributors
 *
 * @date Created: 24th July 2023
 * @date Last Updated: 23th August 2023
 *
 * @version 1.0.0
 *
 * @institute Sapienza University of Rome
 * @cite https://doi.org/10.xxxx/yyyyy
 *
 * @section DEPENDENCIES
 * - Dependency1: Description or version details.
 * - Dependency2: Description or version details.
 *
 * @section LICENSE
 * This file is part of the Aeneas HyperCompute Platform.
 *
 * Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 *
 * @section CHANGELOG
 * @version 1.0.0-dev - 23th August 2023
 * - Initial release
 *
 * @todo
 * - Complete level vector generator function
 * - Add training
 *
 * @see
 * -
 * -
 * -
 *
 */

module class_hvec_gen #(parameter int DI_PARALLEL_W_BITS = 64) (
  input logic [2:0] frame_id,
  input logic [1:0] frame_index,
  output logic [DI_PARALLEL_W_BITS-1:0] class_vec_out
);
  always_comb begin
    case (frame_id)
      0:
        case (frame_index)
          0:
            class_vec_out = 64'b-1077487-1245-1245-1137-1245-1223-124512451003-122112451245-12451245-345-445-12451245-120712451245124511811245-12451245-1245-1245-12456331245-1211943124510711245-1245124512451245-124581-951245-12451245-12011245-1245251-1189-899124564912451245-555853-1039-1245-1105-1245-185;
          1:
            class_vec_out = 64'b-22397-223-223-135-223-217-223223217-223221223-223223127-163-223223-219223223223219223-223223-223-223-223183223-21371223215223-223223223223-223-163-85223-223223-195223-223115-2133922391223223-39201-217-223-187-22321;
          2:
            class_vec_out = 64'b-124-36-126-126-64-126-126-126126114-86126126-126126812-126126-12612612612660126-126126-126-126-12694126-589212644126-126126126126-126-76-66126-126126-116126-12668-118141262412612642100-6-1266-126-44;
        endcase
      1:
        case (frame_index)
          0:
            class_vec_out = 64'b-12455531245-124512451219447-11-113137113912458231245705-1177-1245-34312451215104112431245-823-114179312451245124511792331245197889-11751245-12451245-124575511239751245-1245721-1245124512452372091187-1245-1245-1245-12451245-1245-1245124512451245-1245-12451243;
          1:
            class_vec_out = 64'b-223195223-223223215-51-53-16316119322317922357-219-223-77223215111223223-111-21720122322322322119122319195-217223-223223-223187201211223-22383-2232232231735215-223-223-223-223223-223-223223223223-223-223223;
          2:
            class_vec_out = 64'b-12654126-126126108-76-106-82-26116126-812684-92-126-1061269270118126-16-4258126126126108441266234-88126-126126-1261246642126-126-6-126126126-2218122-126-126-126-126126-126-126126126126-126-126126;
        endcase
      2:
        case (frame_index)
          0:
            class_vec_out = 64'b-1245-8911245124512451245124512451245-1245-1245-1245124512391245731245-124517-1139-1221124512451312451245-72910491245-124512451245-12459251245-1245-11911205-10551241991-1245-12458551245-10912451245-124512458891245-1245-1245-863-1245-124512411245-12451245124512451001;
          1:
            class_vec_out = 64'b-223-189223223223223223223223-223-223-223223221223137223-223-41-217-211223223157223223-179175223-223223223-223199223-223-219211-169219217-223-22323223-163223223-223223207223-223-223-159-223-223223223-223223223223211;
          2:
            class_vec_out = 64'b-1260126126126126126126126-126-126-12612612012644126-126-58-68-11812612628126126-72106126-126126126-126-14126-126-94921612680-126-126-4012624126126-126126120126-126-126-42-126-12698126-12612612612684;
        endcase
      3:
        case (frame_index)
          0:
            class_vec_out = 64'b-12451221-12451245-124571237245-1245-12453321112457571099-12459971245-623-6437331245-12455471063-1245815-12451245-5411245-1219-121312451245-1175-1493031245-1245-1219-1245785-1245-1145-9431245-599211245-12451245-1245-12391239-12451245721823-22745582510711245;
          1:
            class_vec_out = 64'b-223219-223223-223117223-165-223-2231130223-99167-223-2722327-83163223-223195185-223211-223223-97223-219-219223223-159315223-223-223-22351-223-129-189223-7-11223-223223-223-213209-223223-49155121-17211115223;
          2:
            class_vec_out = 64'b-12690-126126-126-485232-126-1263012126-34112-12618126-322484126-12610474-12692-126126-36126-116-110126126-84-5654126-126-122-12652-126-60-56126-2432126-126126-126-86110-1261261090-62496108126;
        endcase
      4:
        case (frame_index)
          0:
            class_vec_out = 64'b1245129357124512411245-1245124512451071-1245-1245-1245-12451245203431-1105-1245-1245-12451245-991-195-227124511718771245-1245-1245-97789-124512451245-11931245141-12453511245-1245-1245-1245124512151229-1245-1245-1245-1245-124562112451245-1233-124596912451245105112451245;
          1:
            class_vec_out = 64'b221-3717223219223-223223223177-223-223-223-22322337-15-193-223-223-223223-215-85-21223209171223-223-223-207-5-223223223-183223181-223-189223-223-223-223223209221-223-223-223-223-223119223223-223-22391223223191223223;
          2:
            class_vec_out = 64'b12636-16126126126-12612612624-126-126-126-126126-3472-100-126-126-126126-92-84-401269098126-126-126-8640-126126126-116126-2-126-22126-126-126-126126120126-126-126-126-126-12638126126-126-12698126126-10126126;
        endcase
      5:
        case (frame_index)
          0:
            class_vec_out = 64'b233-12452311245-1245551-1245785-29-12451245277-1237-12451245-10271245-729-121712451245-1231-7531111193-315-1245881-9751245-1245207-667-12459411245-124512451245124512451245-124512451245-1061-12451245145-1245-1095185-12451245124512451105-1245-12251931245-1245-9091245;
          1:
            class_vec_out = 64'b103-223143223-223-97-223199179-22322333-221-223223-57223-217-219223223-219-179143219-55-223147-209223-223127-111-223123223-223223223223223223-223223223-171-223223115-223-209-55-223223223223169-223-219-87223-223-203223;
          2:
            class_vec_out = 64'b6-12644126-12630-1264814-12612664-104-126126-50126-102-126126126-118261122-12622-100126-1260-74-126108126-126126126126126126-126126126-104-126126-4-126-118-50-12612612012678-126-8444126-126-40126;
        endcase
      6:
        case (frame_index)
          0:
            class_vec_out = 64'b1245-1245-95912451431245-1243-471791115-1245-7791531245-1245-12451207-12431551245-1157-1197-1245-12451087641-1245-124512451245-8551171419-10571245-115512411245-1245-12451245-1245-1245-1245987-46712452856831245-9011235-1245-1245-1245-809116312451245-1231-12451245-477-961;
          1:
            class_vec_out = 64'b223-223-151223-33223-223-737209-223-201115223-223-223223-211-27223-143-221-223-22397183-223-223223223-1332193-187223-215223223-223-223223-223-223-223213-189223-11169223-193211-223-223-223-215201223223-217-223223-49-161;
          2:
            class_vec_out = 64'b126-126-2412666126-126-583054-126-8690126-126-126122-10458126-36-72-126-1269074-126-126126126-8210028126-126100126-126-122126-126-126-12634-141268110126-120116-126-126-126-98104126126-108-126126-82-72;
        endcase
      7:
        case (frame_index)
          0:
            class_vec_out = 64'b1245487-9551245-1245-124579-1245-71-1531245-8871243-1245-12451245-1245-457-83112451239-123112451245437-1245-1245-193-1245-4371245577-767-787743-1245-81-1245-1245115919-12215431245-12455691241124512452851245-12451245-11796531241-1199-579-124591-12451245-1097-1245;
          1:
            class_vec_out = 64'b223127-207223-223-223-185-2231733223-201223-223-223223-22313-57223223-217223223-57-223-223-51-223-113223211107-17357-223-55-223-223211-79-205177223-223-91223223223-19223-223223-179177223-185-189-223161-223223-169-223;
          2:
            class_vec_out = 64'b126100-40126-126-126-90-1263054126-40126-126-126126-126-94-106126126-11412612646-126-126-52-126-11012648-242090-12634-126-12612636-104-18126-1263612612612644126-126126-6612126-98-14-126-16-126126-92-126;
        endcase
    endcase
  end
endmodule