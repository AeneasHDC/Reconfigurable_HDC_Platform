/**
 * @file level_hvec_gen_hdl.hpp
 * @brief This script generates HDL code for generating high-dimensional LEVEL vectors.
 * It is a novel method; for more information, please refer to our paper.
 *
 * @author Saeid Jamili and Marco Angioli
 * @note Author names are listed in alphabetical order.
 * @email <saeid.jamili@uniroma1.it>
 * @email <marco.angioli@uniroma1.it>
 *
 * @contributors
 *
 * @date Created: 24th July 2023
 * @date Last Updated: 23th August 2023
 *
 * @version 1.0.0
 *
 * @institute Sapienza University of Rome
 * @cite https://doi.org/10.xxxx/yyyyy
 *
 * @section DEPENDENCIES
 * - Dependency1: Description or version details.
 * - Dependency2: Description or version details.
 *
 * @section LICENSE
 * This file is part of the Aeneas HyperCompute Platform.
 *
 * Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 *
 * @section CHANGELOG
 * @version 1.0.0-dev - 23th August 2023
 * - Initial release
 *
 * @todo
 * - Complete level vector generator function
 * - Add training
 *
 * @see
 * -
 * -
 * -
 *
 */

module level_hvec_gen #(parameter int DI_PARALLEL_W_BITS = 64) (
  input logic [2:0] frame_index,
  input logic [4:0] frame_id,
  output logic [DI_PARALLEL_W_BITS-1:0] level_vec_out
);
  always_comb begin
    case (frame_index)
      0:
        case (frame_id)
          0:
            level_vec_out = 64'b0001000101000110010001011010001110011011100010011011000100101100;
          1:
            level_vec_out = 64'b0001000101000110010001011010001110011011100010011011000100101100;
          2:
            level_vec_out = 64'b0001000101000110010001011010001110011011100010011011000101101100;
          3:
            level_vec_out = 64'b0001000101000110010001011010001110011011100010011011000101101100;
          4:
            level_vec_out = 64'b0001000101000110010001011010001110011011100010011011000101101100;
          5:
            level_vec_out = 64'b0001000101000110010001011010001110011011100010011011000101101100;
          6:
            level_vec_out = 64'b0001000101000110010001011110001110011011100110011011000101101100;
          7:
            level_vec_out = 64'b0001000101000110010001011110001110011011100110011111000101101100;
          8:
            level_vec_out = 64'b0001010101000110010001011110001110011011100110011111000101101100;
          9:
            level_vec_out = 64'b0001010101000110010001111110001110011011100110011111000101101100;
          10:
            level_vec_out = 64'b0011010101000110010001111110001110011011100110011111000101101100;
          11:
            level_vec_out = 64'b0011110101000110010001111110001110011011100110011111010101101100;
          12:
            level_vec_out = 64'b1011110101000110010011111110101110011011100110011111010101101100;
          13:
            level_vec_out = 64'b1011110101000110010011111110101110011011101110011111010101101100;
          14:
            level_vec_out = 64'b1011110101000110010011111110101110011011101110011111010101101100;
          15:
            level_vec_out = 64'b1011110101000110010011111110101110011011101110011111011101101100;
          16:
            level_vec_out = 64'b1011110101000110010011111110101110011011101110011111011101101100;
          17:
            level_vec_out = 64'b1011110101000110010011111110101110011011101110011111011101101100;
          18:
            level_vec_out = 64'b1011111101010110010011111110101110011011111110011111011101101100;
          19:
            level_vec_out = 64'b1011111101010110010011111110111110011011111111011111111101101100;
          20:
            level_vec_out = 64'b1011111101010110010011111110111111011011111111011111111101101110;
          21:
            level_vec_out = 64'b1011111101010110010011111110111111011011111111011111111101101110;
          22:
            level_vec_out = 64'b1011111101010110010111111111111111011011111111011111111111101110;
          23:
            level_vec_out = 64'b1011111101010110010111111111111111011011111111011111111111101110;
          24:
            level_vec_out = 64'b1011111101110110010111111111111111011011111111011111111111101110;
          25:
            level_vec_out = 64'b1011111111110110111111111111111111011111111111011111111111101110;
          26:
            level_vec_out = 64'b1011111111111110111111111111111111011111111111011111111111101110;
          27:
            level_vec_out = 64'b1011111111111110111111111111111111011111111111011111111111101111;
          28:
            level_vec_out = 64'b1011111111111110111111111111111111111111111111011111111111101111;
          29:
            level_vec_out = 64'b1011111111111110111111111111111111111111111111011111111111101111;
          30:
            level_vec_out = 64'b1111111111111110111111111111111111111111111111111111111111111111;
          31:
            level_vec_out = 64'b1111111111111110111111111111111111111111111111111111111111111111;
        endcase
      1:
        case (frame_id)
          0:
            level_vec_out = 64'b0111000000100110000111011100111011001011101110101001011111000110;
          1:
            level_vec_out = 64'b0111000000100110000111011101111011001011101110101001011111000110;
          2:
            level_vec_out = 64'b0111000000100110000111011101111011001011111110101001011111000110;
          3:
            level_vec_out = 64'b0111000000100110000111011101111011001011111111101001011111000110;
          4:
            level_vec_out = 64'b0111000000100110000111011101111011001011111111101011011111000111;
          5:
            level_vec_out = 64'b0111000000100110000111011101111011001011111111101011011111000111;
          6:
            level_vec_out = 64'b0111000001100110000111011101111011001011111111101011011111000111;
          7:
            level_vec_out = 64'b0111000001100110000111011101111011001011111111101111011111000111;
          8:
            level_vec_out = 64'b0111000001100111000111011101111011001011111111101111011111000111;
          9:
            level_vec_out = 64'b1111000001101111000111011101111011001011111111101111011111000111;
          10:
            level_vec_out = 64'b1111000011101111000111011101111011001011111111101111011111000111;
          11:
            level_vec_out = 64'b1111000011101111000111011101111011001011111111101111011111000111;
          12:
            level_vec_out = 64'b1111000011101111000111011101111011001011111111101111011111000111;
          13:
            level_vec_out = 64'b1111000011101111000111011101111011001011111111101111011111000111;
          14:
            level_vec_out = 64'b1111000011101111000111011101111111001011111111101111011111000111;
          15:
            level_vec_out = 64'b1111001011101111000111011101111111001011111111101111011111000111;
          16:
            level_vec_out = 64'b1111001111101111100111011111111111001011111111101111011111000111;
          17:
            level_vec_out = 64'b1111001111101111100111011111111111001111111111101111011111100111;
          18:
            level_vec_out = 64'b1111001111101111100111011111111111001111111111101111011111100111;
          19:
            level_vec_out = 64'b1111011111101111110111011111111111001111111111101111011111100111;
          20:
            level_vec_out = 64'b1111011111101111110111011111111111011111111111101111011111100111;
          21:
            level_vec_out = 64'b1111011111101111111111011111111111011111111111111111011111100111;
          22:
            level_vec_out = 64'b1111011111111111111111011111111111011111111111111111011111100111;
          23:
            level_vec_out = 64'b1111011111111111111111011111111111011111111111111111111111100111;
          24:
            level_vec_out = 64'b1111011111111111111111011111111111011111111111111111111111100111;
          25:
            level_vec_out = 64'b1111011111111111111111011111111111011111111111111111111111110111;
          26:
            level_vec_out = 64'b1111011111111111111111011111111111011111111111111111111111110111;
          27:
            level_vec_out = 64'b1111011111111111111111111111111111011111111111111111111111110111;
          28:
            level_vec_out = 64'b1111011111111111111111111111111111011111111111111111111111111111;
          29:
            level_vec_out = 64'b1111111111111111111111111111111111011111111111111111111111111111;
          30:
            level_vec_out = 64'b1111111111111111111111111111111111011111111111111111111111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111011111111111111111111111111111;
        endcase
      2:
        case (frame_id)
          0:
            level_vec_out = 64'b0110011011111111100011110001100111100001101110111011001110111010;
          1:
            level_vec_out = 64'b0110011011111111100011110001100111100001101110111011001110111010;
          2:
            level_vec_out = 64'b0110011011111111100011110101100111100001101110111011001110111010;
          3:
            level_vec_out = 64'b0110011011111111100011110101100111100001111110111011001110111010;
          4:
            level_vec_out = 64'b0110011011111111100011110101100111100001111110111011001110111010;
          5:
            level_vec_out = 64'b0110011011111111100011110111100111100001111110111011001110111010;
          6:
            level_vec_out = 64'b0110011011111111100011110111100111100001111110111011001110111110;
          7:
            level_vec_out = 64'b0110111011111111100011110111100111100001111110111011001110111110;
          8:
            level_vec_out = 64'b0110111011111111100011111111100111100001111110111011001110111110;
          9:
            level_vec_out = 64'b0110111011111111100011111111110111100001111110111011001110111110;
          10:
            level_vec_out = 64'b0110111011111111100011111111110111100101111110111011001111111110;
          11:
            level_vec_out = 64'b0110111011111111100011111111110111100101111110111011011111111110;
          12:
            level_vec_out = 64'b0110111011111111100011111111110111100101111110111011011111111110;
          13:
            level_vec_out = 64'b0110111011111111100011111111110111100101111110111011011111111110;
          14:
            level_vec_out = 64'b0110111011111111110011111111110111100101111110111011011111111110;
          15:
            level_vec_out = 64'b0110111111111111111011111111110111100101111110111011011111111110;
          16:
            level_vec_out = 64'b0110111111111111111011111111110111100101111110111011011111111110;
          17:
            level_vec_out = 64'b0110111111111111111011111111110111100101111110111011011111111110;
          18:
            level_vec_out = 64'b0110111111111111111011111111110111100101111110111011011111111110;
          19:
            level_vec_out = 64'b0110111111111111111011111111110111100101111110111011011111111110;
          20:
            level_vec_out = 64'b0110111111111111111011111111110111101101111110111011011111111110;
          21:
            level_vec_out = 64'b0110111111111111111011111111110111101101111110111011011111111110;
          22:
            level_vec_out = 64'b0110111111111111111011111111110111101101111110111011011111111111;
          23:
            level_vec_out = 64'b1110111111111111111011111111110111101101111110111011011111111111;
          24:
            level_vec_out = 64'b1110111111111111111011111111110111111101111110111011011111111111;
          25:
            level_vec_out = 64'b1110111111111111111111111111110111111101111110111011011111111111;
          26:
            level_vec_out = 64'b1110111111111111111111111111111111111101111110111011011111111111;
          27:
            level_vec_out = 64'b1110111111111111111111111111111111111101111111111111011111111111;
          28:
            level_vec_out = 64'b1110111111111111111111111111111111111101111111111111011111111111;
          29:
            level_vec_out = 64'b1110111111111111111111111111111111111101111111111111011111111111;
          30:
            level_vec_out = 64'b1110111111111111111111111111111111111101111111111111011111111111;
          31:
            level_vec_out = 64'b1110111111111111111111111111111111111111111111111111111111111111;
        endcase
      3:
        case (frame_id)
          0:
            level_vec_out = 64'b1100101111100000101011110110010001101000110000000011000111110001;
          1:
            level_vec_out = 64'b1110101111100000101011110110010001101000110000000011000111110001;
          2:
            level_vec_out = 64'b1110101111100000101011110110010001101000110100000011000111110001;
          3:
            level_vec_out = 64'b1111101111100000101011110110010001101000110100000111000111110011;
          4:
            level_vec_out = 64'b1111101111100000101011110110110001101000110100010111000111110011;
          5:
            level_vec_out = 64'b1111101111100100101011110110110001101000110101010111000111110011;
          6:
            level_vec_out = 64'b1111101111100100101011110110110001111000110101010111000111110011;
          7:
            level_vec_out = 64'b1111101111100100101011110110110001111000110101110111000111110011;
          8:
            level_vec_out = 64'b1111101111100100101111111110110001111000110101110111000111110011;
          9:
            level_vec_out = 64'b1111101111100100101111111110110001111000110101111111000111110011;
          10:
            level_vec_out = 64'b1111101111100100101111111111110001111000110101111111001111110011;
          11:
            level_vec_out = 64'b1111101111110100101111111111110001111000110101111111001111110011;
          12:
            level_vec_out = 64'b1111101111110100101111111111110001111000110111111111001111110011;
          13:
            level_vec_out = 64'b1111101111110100101111111111110001111001110111111111001111110011;
          14:
            level_vec_out = 64'b1111101111110110101111111111110001111001110111111111001111110011;
          15:
            level_vec_out = 64'b1111101111110110101111111111110001111001110111111111001111110011;
          16:
            level_vec_out = 64'b1111101111110110101111111111110001111001110111111111001111110011;
          17:
            level_vec_out = 64'b1111101111110110101111111111110001111001110111111111001111110011;
          18:
            level_vec_out = 64'b1111101111110110101111111111110101111001110111111111001111110011;
          19:
            level_vec_out = 64'b1111101111110110101111111111110101111001110111111111001111110011;
          20:
            level_vec_out = 64'b1111101111110110101111111111110101111001110111111111001111110011;
          21:
            level_vec_out = 64'b1111101111110110101111111111110101111001110111111111001111110011;
          22:
            level_vec_out = 64'b1111101111110110111111111111111101111001110111111111001111110011;
          23:
            level_vec_out = 64'b1111101111111110111111111111111101111001110111111111001111110011;
          24:
            level_vec_out = 64'b1111101111111110111111111111111101111001110111111111011111110111;
          25:
            level_vec_out = 64'b1111101111111110111111111111111101111001110111111111011111110111;
          26:
            level_vec_out = 64'b1111101111111110111111111111111101111011110111111111011111111111;
          27:
            level_vec_out = 64'b1111101111111110111111111111111101111011110111111111011111111111;
          28:
            level_vec_out = 64'b1111111111111110111111111111111101111011110111111111011111111111;
          29:
            level_vec_out = 64'b1111111111111111111111111111111101111011110111111111111111111111;
          30:
            level_vec_out = 64'b1111111111111111111111111111111101111011110111111111111111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111101111111111111111111111111111111;
        endcase
      4:
        case (frame_id)
          0:
            level_vec_out = 64'b0001110111100001011100101100010000011010001000001000001000111100;
          1:
            level_vec_out = 64'b0001110111100001011100101100010000011111001000001000001100111100;
          2:
            level_vec_out = 64'b0001110111100001011100101100110000011111001000001000001100111100;
          3:
            level_vec_out = 64'b0001110111100001111100101100110000011111001000001000001100111100;
          4:
            level_vec_out = 64'b0001110111100001111100101100110000011111001100001001001100111100;
          5:
            level_vec_out = 64'b0001110111100001111100101100110000011111001110011001001100111100;
          6:
            level_vec_out = 64'b0001110111100001111100101100111000011111001110011001011100111100;
          7:
            level_vec_out = 64'b0001110111100001111100101100111000011111001110011001111100111100;
          8:
            level_vec_out = 64'b0001110111100001111100101100111000011111001110011001111100111100;
          9:
            level_vec_out = 64'b0001110111100001111100101100111000011111001110011001111100111100;
          10:
            level_vec_out = 64'b0001110111100001111100101100111000011111001110011001111100111100;
          11:
            level_vec_out = 64'b0001110111100001111100101100111000011111001110011011111100111110;
          12:
            level_vec_out = 64'b0001111111100001111100101100111000111111001110011011111100111111;
          13:
            level_vec_out = 64'b0001111111100001111110101100111000111111001110011011111100111111;
          14:
            level_vec_out = 64'b0001111111100001111110101100111000111111001110011011111100111111;
          15:
            level_vec_out = 64'b0001111111100001111110101100111000111111001110111011111100111111;
          16:
            level_vec_out = 64'b0001111111100001111110101100111001111111011110111011111100111111;
          17:
            level_vec_out = 64'b0001111111100001111111111100111001111111011110111011111100111111;
          18:
            level_vec_out = 64'b0001111111100001111111111100111001111111011110111011111100111111;
          19:
            level_vec_out = 64'b0001111111100001111111111100111001111111011110111011111100111111;
          20:
            level_vec_out = 64'b0001111111100101111111111100111001111111011110111011111100111111;
          21:
            level_vec_out = 64'b0011111111110101111111111101111001111111011110111111111100111111;
          22:
            level_vec_out = 64'b0011111111110101111111111101111001111111011110111111111100111111;
          23:
            level_vec_out = 64'b0011111111110111111111111101111001111111011110111111111100111111;
          24:
            level_vec_out = 64'b0011111111110111111111111101111101111111011110111111111100111111;
          25:
            level_vec_out = 64'b0011111111110111111111111101111101111111011110111111111100111111;
          26:
            level_vec_out = 64'b0011111111110111111111111101111101111111011110111111111100111111;
          27:
            level_vec_out = 64'b0011111111110111111111111101111101111111011110111111111110111111;
          28:
            level_vec_out = 64'b0011111111110111111111111101111101111111011111111111111110111111;
          29:
            level_vec_out = 64'b0111111111110111111111111101111101111111011111111111111110111111;
          30:
            level_vec_out = 64'b1111111111110111111111111101111101111111011111111111111111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111101111111011111111111111111111111;
        endcase
      5:
        case (frame_id)
          0:
            level_vec_out = 64'b0001100101001100101000000000111001100010000110110011101110001011;
          1:
            level_vec_out = 64'b0001100101001110101000000000111001100010000110110011111110001011;
          2:
            level_vec_out = 64'b1001101101001110101000000000111001100010000110110011111110001011;
          3:
            level_vec_out = 64'b1001101101001110101000000000111001100010000110110011111110001011;
          4:
            level_vec_out = 64'b1001101101001110101000000010111001100010000110110011111110001011;
          5:
            level_vec_out = 64'b1001101101001110101000010010111001100010000110110011111110101011;
          6:
            level_vec_out = 64'b1001101101001110101000010010111001100010000110111011111110101011;
          7:
            level_vec_out = 64'b1001101101001110111000010010111001100010000110111011111110101011;
          8:
            level_vec_out = 64'b1001101101001110111000010010111001100010000110111011111110101011;
          9:
            level_vec_out = 64'b1001101101001110111000010010111001100010000110111011111110101011;
          10:
            level_vec_out = 64'b1001101101011110111000010010111001100010000110111011111110101011;
          11:
            level_vec_out = 64'b1001101101011110111000010010111001100010010110111011111110101011;
          12:
            level_vec_out = 64'b1001101101011110111000010010111001100010010110111011111110101011;
          13:
            level_vec_out = 64'b1001101101011110111001010010111001100010010110111011111110101111;
          14:
            level_vec_out = 64'b1001101101011110111001011010111001100110010110111011111110101111;
          15:
            level_vec_out = 64'b1001101101011111111001011010111001100110010110111011111110101111;
          16:
            level_vec_out = 64'b1001101101011111111001011010111001100110010111111011111110101111;
          17:
            level_vec_out = 64'b1001101101011111111001011010111001100111010111111111111110101111;
          18:
            level_vec_out = 64'b1011101101011111111001011010111101100111010111111111111110101111;
          19:
            level_vec_out = 64'b1011101101011111111011011010111101100111010111111111111110101111;
          20:
            level_vec_out = 64'b1011101101011111111011011010111101100111110111111111111110101111;
          21:
            level_vec_out = 64'b1011101101011111111011011010111101100111110111111111111110101111;
          22:
            level_vec_out = 64'b1011101101011111111011011010111101100111110111111111111110101111;
          23:
            level_vec_out = 64'b1011101101011111111111111010111101101111110111111111111111101111;
          24:
            level_vec_out = 64'b1011101101011111111111111110111101101111111111111111111111101111;
          25:
            level_vec_out = 64'b1011101101011111111111111110111101101111111111111111111111101111;
          26:
            level_vec_out = 64'b1011101101011111111111111110111101111111111111111111111111101111;
          27:
            level_vec_out = 64'b1011101101011111111111111110111101111111111111111111111111101111;
          28:
            level_vec_out = 64'b1011111101011111111111111110111101111111111111111111111111111111;
          29:
            level_vec_out = 64'b1011111111011111111111111110111101111111111111111111111111111111;
          30:
            level_vec_out = 64'b1111111111011111111111111110111101111111111111111111111111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111101111111111111111111111111111111;
        endcase
      6:
        case (frame_id)
          0:
            level_vec_out = 64'b0010010101100101010110110110111011000111010011000111101010011111;
          1:
            level_vec_out = 64'b0011010101100101010110110110111011000111010011000111101010011111;
          2:
            level_vec_out = 64'b0011010101100101010110110111111011000111010011000111101010011111;
          3:
            level_vec_out = 64'b0011010101100101010110110111111011000111011011000111101010011111;
          4:
            level_vec_out = 64'b0011010101100111010110110111111011000111011011000111101010011111;
          5:
            level_vec_out = 64'b0011010101100111010110110111111011000111011011000111101010011111;
          6:
            level_vec_out = 64'b0011010101100111010110110111111011000111011011000111101010011111;
          7:
            level_vec_out = 64'b0011010101100111010110110111111011000111011011000111101010011111;
          8:
            level_vec_out = 64'b0011010101100111010110110111111011000111011011000111101010111111;
          9:
            level_vec_out = 64'b0011010101100111011110110111111011000111011011000111101010111111;
          10:
            level_vec_out = 64'b0011010101100111011110110111111011000111011011000111101110111111;
          11:
            level_vec_out = 64'b0011010101100111011110110111111011000111011011010111101110111111;
          12:
            level_vec_out = 64'b0011010101100111011110110111111011000111011011010111101110111111;
          13:
            level_vec_out = 64'b0111110101100111011110110111111011000111011011010111111110111111;
          14:
            level_vec_out = 64'b0111110101100111011110110111111011100111011111010111111110111111;
          15:
            level_vec_out = 64'b1111110101100111011110110111111011100111011111010111111110111111;
          16:
            level_vec_out = 64'b1111110101100111011110110111111011110111011111010111111110111111;
          17:
            level_vec_out = 64'b1111110101100111011110110111111011110111111111010111111110111111;
          18:
            level_vec_out = 64'b1111111101100111011110111111111011110111111111010111111110111111;
          19:
            level_vec_out = 64'b1111111101100111011110111111111111110111111111010111111110111111;
          20:
            level_vec_out = 64'b1111111101100111011110111111111111111111111111010111111111111111;
          21:
            level_vec_out = 64'b1111111101100111011110111111111111111111111111010111111111111111;
          22:
            level_vec_out = 64'b1111111101100111011110111111111111111111111111010111111111111111;
          23:
            level_vec_out = 64'b1111111101100111011110111111111111111111111111010111111111111111;
          24:
            level_vec_out = 64'b1111111101100111011110111111111111111111111111010111111111111111;
          25:
            level_vec_out = 64'b1111111101100111011110111111111111111111111111010111111111111111;
          26:
            level_vec_out = 64'b1111111101100111011110111111111111111111111111111111111111111111;
          27:
            level_vec_out = 64'b1111111111110111111110111111111111111111111111111111111111111111;
          28:
            level_vec_out = 64'b1111111111110111111110111111111111111111111111111111111111111111;
          29:
            level_vec_out = 64'b1111111111111111111110111111111111111111111111111111111111111111;
          30:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        endcase
      7:
        case (frame_id)
          0:
            level_vec_out = 64'b1011001011011010111010010011111011000110111001111110110011000100;
          1:
            level_vec_out = 64'b1011001011011010111010010011111011000110111001111110110011000100;
          2:
            level_vec_out = 64'b1011001011011010111010010011111011000110111001111110110011000100;
          3:
            level_vec_out = 64'b1011001011111010111010010011111011000110111001111110110011000100;
          4:
            level_vec_out = 64'b1011001011111010111010010011111011000110111001111110110011000100;
          5:
            level_vec_out = 64'b1011001011111010111010110011111011000110111001111110110011000100;
          6:
            level_vec_out = 64'b1011001011111010111010110011111011000110111001111110110011000100;
          7:
            level_vec_out = 64'b1011001111111010111011110011111011000110111001111110110011000100;
          8:
            level_vec_out = 64'b1011001111111011111011110011111011000110111011111110110011000100;
          9:
            level_vec_out = 64'b1011001111111011111011110011111111000110111011111111110011000100;
          10:
            level_vec_out = 64'b1011001111111011111011110011111111000110111011111111110011000100;
          11:
            level_vec_out = 64'b1011001111111011111011110011111111000110111011111111110011000100;
          12:
            level_vec_out = 64'b1011001111111011111011110011111111000110111111111111110011000100;
          13:
            level_vec_out = 64'b1011001111111011111011110011111111000110111111111111110011000100;
          14:
            level_vec_out = 64'b1011001111111011111011110011111111000110111111111111110011000101;
          15:
            level_vec_out = 64'b1011001111111011111011110011111111000110111111111111110011100101;
          16:
            level_vec_out = 64'b1011001111111011111011110011111111010110111111111111110011100101;
          17:
            level_vec_out = 64'b1011001111111011111011110011111111010110111111111111111011100101;
          18:
            level_vec_out = 64'b1011001111111011111011110011111111010110111111111111111011100101;
          19:
            level_vec_out = 64'b1011001111111111111011110011111111010110111111111111111011100101;
          20:
            level_vec_out = 64'b1011001111111111111011110011111111010110111111111111111011100101;
          21:
            level_vec_out = 64'b1011001111111111111011111011111111011110111111111111111011100101;
          22:
            level_vec_out = 64'b1011001111111111111011111011111111011111111111111111111011100101;
          23:
            level_vec_out = 64'b1011001111111111111011111011111111011111111111111111111011100101;
          24:
            level_vec_out = 64'b1011001111111111111011111011111111011111111111111111111111100101;
          25:
            level_vec_out = 64'b1011001111111111111011111111111111111111111111111111111111100101;
          26:
            level_vec_out = 64'b1011001111111111111111111111111111111111111111111111111111100101;
          27:
            level_vec_out = 64'b1011001111111111111111111111111111111111111111111111111111100101;
          28:
            level_vec_out = 64'b1111001111111111111111111111111111111111111111111111111111110101;
          29:
            level_vec_out = 64'b1111011111111111111111111111111111111111111111111111111111111101;
          30:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111101;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111101;
        endcase
    endcase
  end
endmodule