----
 -- @file level_hvec_gen_hdl.hpp
 -- @brief This script generates HDL code for generating high-dimensional LEVEL vectors.
 -- It is a novel method; for more information, please refer to our paper.
 --
 -- @author Saeid Jamili and Marco Angioli
 -- @note Author names are listed in alphabetical order.
 -- @email <saeid.jamili@uniroma1.it>
 -- @email <marco.angioli@uniroma1.it>
 --
 -- @contributors
 --
 -- @date Created: 24th July 2023
 -- @date Last Updated: 23th August 2023
 --
 -- @version 1.0.0
 --
 -- @institute Sapienza University of Rome
 -- @cite https://doi.org/10.xxxx/yyyyy
 --
 -- @section DEPENDENCIES
 -- - Dependency1: Description or version details.
 -- - Dependency2: Description or version details.
 --
 -- @section LICENSE
 -- This file is part of the Aeneas HyperCompute Platform.
 --
 -- Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 --
 -- @section CHANGELOG
 -- @version 1.0.0-dev - 23th August 2023
 -- - Initial release
 --
 -- @todo
 -- - Complete level vector generator function
 -- - Add training
 --
 -- @see
 -- -
 -- -
 -- -
 --
 --

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity level_vec_gen is
    Port ( level_vec_out : out  STD_LOGIC_VECTOR (63 downto 0);
           frame_index : in  STD_LOGIC_VECTOR (2 downto 0);
           frame_id : in  STD_LOGIC_VECTOR (4 downto 0));
end level_vec_gen;

architecture Behavioral of level_vec_gen is
begin
    process (frame_index, frame_id)
    begin
        -- Update this function to match your requirements
        case frame_index is
            when "000" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1000100110001011101101101111001110000110111001011001010000010000";
                    when "00001" => level_vec_out <= "1000100110001011101101101111001110000110111001011001010000010001";
                    when "00010" => level_vec_out <= "1000100110001011101101101111001110000110111001011001010000010001";
                    when "00011" => level_vec_out <= "1000100111001011101111101111011111000110111001011001010000010011";
                    when "00100" => level_vec_out <= "1000100111001011101111101111011111000110111001011001010000010011";
                    when "00101" => level_vec_out <= "1000100111001011101111101111011111000110111101011001010000010011";
                    when "00110" => level_vec_out <= "1000100111001011101111111111011111000110111101011001010000010011";
                    when "00111" => level_vec_out <= "1010100111001011101111111111011111000110111101011001010000010011";
                    when "01000" => level_vec_out <= "1010100111001011101111111111011111000111111101011001010000010011";
                    when "01001" => level_vec_out <= "1011100111001011101111111111011111000111111101011001010000010011";
                    when "01010" => level_vec_out <= "1011100111001011101111111111011111000111111101011001010000011011";
                    when "01011" => level_vec_out <= "1011100111001011101111111111011111000111111101011001010000011011";
                    when "01100" => level_vec_out <= "1011100111001011101111111111011111000111111101011001010100011011";
                    when "01101" => level_vec_out <= "1011100111001011101111111111011111000111111101011001010100111011";
                    when "01110" => level_vec_out <= "1011100111001011101111111111011111000111111101111001010100111111";
                    when "01111" => level_vec_out <= "1011100111001011101111111111011111010111111101111001010110111111";
                    when "10000" => level_vec_out <= "1011100111001011101111111111011111010111111101111001010110111111";
                    when "10001" => level_vec_out <= "1011100111001011101111111111011111010111111101111001010111111111";
                    when "10010" => level_vec_out <= "1011100111001011101111111111011111010111111101111001110111111111";
                    when "10011" => level_vec_out <= "1011100111001011101111111111011111011111111111111011110111111111";
                    when "10100" => level_vec_out <= "1011100111001011101111111111011111011111111111111011110111111111";
                    when "10101" => level_vec_out <= "1011100111001011111111111111011111011111111111111011110111111111";
                    when "10110" => level_vec_out <= "1011100111001011111111111111011111011111111111111011110111111111";
                    when "10111" => level_vec_out <= "1011100111001011111111111111011111011111111111111011111111111111";
                    when "11000" => level_vec_out <= "1111100111001011111111111111011111011111111111111011111111111111";
                    when "11001" => level_vec_out <= "1111100111001011111111111111011111111111111111111011111111111111";
                    when "11010" => level_vec_out <= "1111100111001011111111111111011111111111111111111011111111111111";
                    when "11011" => level_vec_out <= "1111100111001011111111111111011111111111111111111011111111111111";
                    when "11100" => level_vec_out <= "1111100111101111111111111111011111111111111111111011111111111111";
                    when "11101" => level_vec_out <= "1111100111101111111111111111011111111111111111111011111111111111";
                    when "11110" => level_vec_out <= "1111110111101111111111111111011111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111110111101111111111111111011111111111111111111111111111111111";
                when others => null;
                end case;
            when "001" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1001010001110010001111001010001010011001110111111001100100101110";
                    when "00001" => level_vec_out <= "1001010001110010001111001010001010011101110111111001100100101110";
                    when "00010" => level_vec_out <= "1011010001110010001111001010001010011101110111111001100110101110";
                    when "00011" => level_vec_out <= "1011010001110010001111001010001010011101110111111001100110101110";
                    when "00100" => level_vec_out <= "1111010011110010001111001010001010011101110111111001100110101110";
                    when "00101" => level_vec_out <= "1111010011110010001111001010001010011101110111111001100110101110";
                    when "00110" => level_vec_out <= "1111010011110010001111001010001010011101110111111001101110101110";
                    when "00111" => level_vec_out <= "1111010011110110001111001010001010011101110111111011101110101110";
                    when "01000" => level_vec_out <= "1111110011110110001111001010001010011101110111111011111110101110";
                    when "01001" => level_vec_out <= "1111110011110110001111001010001010011101110111111011111110101110";
                    when "01010" => level_vec_out <= "1111111011111110001111001010001010011101110111111011111110101111";
                    when "01011" => level_vec_out <= "1111111011111110001111001010001011011101110111111011111110101111";
                    when "01100" => level_vec_out <= "1111111011111110001111001010001011011101110111111011111110101111";
                    when "01101" => level_vec_out <= "1111111011111110001111001010001011011101110111111011111110101111";
                    when "01110" => level_vec_out <= "1111111011111110001111001010001011011101110111111011111110101111";
                    when "01111" => level_vec_out <= "1111111011111110001111001010001011011101110111111011111110101111";
                    when "10000" => level_vec_out <= "1111111011111110101111001010101011011101110111111011111110101111";
                    when "10001" => level_vec_out <= "1111111011111110101111001010101011011101111111111011111110101111";
                    when "10010" => level_vec_out <= "1111111011111110101111001011101011011101111111111011111110111111";
                    when "10011" => level_vec_out <= "1111111011111110101111001111101011011101111111111011111110111111";
                    when "10100" => level_vec_out <= "1111111011111110101111001111101011011101111111111011111110111111";
                    when "10101" => level_vec_out <= "1111111011111110101111001111101011011101111111111011111111111111";
                    when "10110" => level_vec_out <= "1111111011111110101111001111101011011101111111111011111111111111";
                    when "10111" => level_vec_out <= "1111111011111110101111001111101111011101111111111111111111111111";
                    when "11000" => level_vec_out <= "1111111011111110101111001111101111011101111111111111111111111111";
                    when "11001" => level_vec_out <= "1111111011111110111111001111101111011101111111111111111111111111";
                    when "11010" => level_vec_out <= "1111111111111110111111001111101111111101111111111111111111111111";
                    when "11011" => level_vec_out <= "1111111111111110111111001111101111111101111111111111111111111111";
                    when "11100" => level_vec_out <= "1111111111111110111111001111101111111111111111111111111111111111";
                    when "11101" => level_vec_out <= "1111111111111111111111011111101111111111111111111111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "010" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1010010100010001111000110101111101111010011101010111000011100010";
                    when "00001" => level_vec_out <= "1010010100010001111000110101111101111110011101010111000011100010";
                    when "00010" => level_vec_out <= "1010010100010001111000110101111101111110011101010111000011100010";
                    when "00011" => level_vec_out <= "1010010100010001111000110101111101111110011101010111000011100010";
                    when "00100" => level_vec_out <= "1010010100010001111000110101111101111110011101010111000011100010";
                    when "00101" => level_vec_out <= "1010110100010001111000110101111101111110011101010111100011100010";
                    when "00110" => level_vec_out <= "1010110100010001111000110101111101111110011101010111100011100010";
                    when "00111" => level_vec_out <= "1010110100010001111100110101111101111110011101010111110011100010";
                    when "01000" => level_vec_out <= "1010110100010001111100110101111101111110011101010111110011100010";
                    when "01001" => level_vec_out <= "1010110100010001111100111101111101111110011101010111110011100010";
                    when "01010" => level_vec_out <= "1010110100011001111100111101111101111110011101010111110011100010";
                    when "01011" => level_vec_out <= "1010110100011001111100111101111101111110011101010111110011100010";
                    when "01100" => level_vec_out <= "1010110100011001111100111101111101111110011101010111110011100010";
                    when "01101" => level_vec_out <= "1110110100011011111100111101111101111110011101010111110011100011";
                    when "01110" => level_vec_out <= "1110111100011011111100111101111101111110011111010111110011100011";
                    when "01111" => level_vec_out <= "1110111100011011111100111101111101111110011111010111110011100011";
                    when "10000" => level_vec_out <= "1110111100011011111100111111111101111110011111010111110011100011";
                    when "10001" => level_vec_out <= "1110111100011011111110111111111101111110011111010111110011100011";
                    when "10010" => level_vec_out <= "1110111100011011111110111111111101111110011111010111110011100011";
                    when "10011" => level_vec_out <= "1111111100011011111110111111111101111110011111010111110011100011";
                    when "10100" => level_vec_out <= "1111111100111011111110111111111101111110011111010111110011100011";
                    when "10101" => level_vec_out <= "1111111100111011111110111111111101111110011111110111110011110011";
                    when "10110" => level_vec_out <= "1111111110111011111110111111111101111110011111110111110011111011";
                    when "10111" => level_vec_out <= "1111111110111011111110111111111101111110011111110111110011111011";
                    when "11000" => level_vec_out <= "1111111110111011111110111111111101111110011111111111111011111011";
                    when "11001" => level_vec_out <= "1111111110111011111110111111111101111110011111111111111011111011";
                    when "11010" => level_vec_out <= "1111111111111011111110111111111111111110011111111111111011111011";
                    when "11011" => level_vec_out <= "1111111111111011111110111111111111111110111111111111111011111011";
                    when "11100" => level_vec_out <= "1111111111111011111110111111111111111110111111111111111011111011";
                    when "11101" => level_vec_out <= "1111111111111011111110111111111111111111111111111111111011111011";
                    when "11110" => level_vec_out <= "1111111111111111111110111111111111111111111111111111111011111011";
                    when "11111" => level_vec_out <= "1111111111111111111110111111111111111111111111111111111011111111";
                when others => null;
                end case;
            when "011" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0011011101000101101101110010011011000001011111001110111010000110";
                    when "00001" => level_vec_out <= "0011011101000101101101110010011011100001011111001110111010000111";
                    when "00010" => level_vec_out <= "0011011101000101101101110010011011100001011111001110111010000111";
                    when "00011" => level_vec_out <= "0011011101000101101101110010011011100001011111011110111010000111";
                    when "00100" => level_vec_out <= "0011011101000101101101110010011011100001011111011110111010000111";
                    when "00101" => level_vec_out <= "0011011101000101101101110010011011101001011111011110111010000111";
                    when "00110" => level_vec_out <= "0011011101000101101101111010011011101001011111011110111010100111";
                    when "00111" => level_vec_out <= "0011011101000101111101111010011011101001011111011110111010100111";
                    when "01000" => level_vec_out <= "0011011101000101111101111010011011101001011111011111111010100111";
                    when "01001" => level_vec_out <= "0011011101001101111101111010111011101001011111011111111010100111";
                    when "01010" => level_vec_out <= "0011011101001101111101111010111011101001011111011111111010100111";
                    when "01011" => level_vec_out <= "0011011101001101111101111010111011101001011111011111111110100111";
                    when "01100" => level_vec_out <= "0011011101001101111101111010111011101001011111011111111110100111";
                    when "01101" => level_vec_out <= "0011011101001101111101111010111011101001011111011111111110101111";
                    when "01110" => level_vec_out <= "0011011101001101111111111010111011101001111111011111111110101111";
                    when "01111" => level_vec_out <= "1011111101011101111111111010111011101001111111011111111110101111";
                    when "10000" => level_vec_out <= "1011111101011101111111111010111011101001111111011111111110101111";
                    when "10001" => level_vec_out <= "1011111101011101111111111010111011101001111111011111111110101111";
                    when "10010" => level_vec_out <= "1111111101011101111111111011111011101001111111011111111110101111";
                    when "10011" => level_vec_out <= "1111111101011101111111111011111011101001111111011111111110101111";
                    when "10100" => level_vec_out <= "1111111101011101111111111011111011101001111111011111111110111111";
                    when "10101" => level_vec_out <= "1111111101011101111111111011111011101001111111011111111110111111";
                    when "10110" => level_vec_out <= "1111111101111101111111111011111011101101111111111111111110111111";
                    when "10111" => level_vec_out <= "1111111101111101111111111011111011101101111111111111111110111111";
                    when "11000" => level_vec_out <= "1111111101111101111111111011111011101101111111111111111110111111";
                    when "11001" => level_vec_out <= "1111111101111101111111111111111011101101111111111111111110111111";
                    when "11010" => level_vec_out <= "1111111101111101111111111111111011101101111111111111111110111111";
                    when "11011" => level_vec_out <= "1111111101111101111111111111111011101101111111111111111110111111";
                    when "11100" => level_vec_out <= "1111111101111101111111111111111111101101111111111111111110111111";
                    when "11101" => level_vec_out <= "1111111111111111111111111111111111101101111111111111111110111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111101101111111111111111110111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111101111111111111111111111111";
                when others => null;
                end case;
            when "100" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0100101100101001010010011000001110111110111001000011111000001010";
                    when "00001" => level_vec_out <= "0100101100101001010010011000001110111110111001100011111000001010";
                    when "00010" => level_vec_out <= "0101101100101001010010011000001110111110111001100011111000001010";
                    when "00011" => level_vec_out <= "0101101100101001010010011000001110111110111001100011111000001010";
                    when "00100" => level_vec_out <= "0101101100101001010010011000001111111110111001100011111000001010";
                    when "00101" => level_vec_out <= "0101101100101001010010011001001111111110111001100011111000001010";
                    when "00110" => level_vec_out <= "0101111100101001010110011001001111111110111001100011111000101010";
                    when "00111" => level_vec_out <= "0101111100101001010110011001001111111110111001100011111000101010";
                    when "01000" => level_vec_out <= "0101111100101001010110011001001111111110111001100011111000101010";
                    when "01001" => level_vec_out <= "0101111100101111010110011001001111111110111001100011111000101010";
                    when "01010" => level_vec_out <= "0101111100101111010110111001001111111110111001100011111000101010";
                    when "01011" => level_vec_out <= "0101111100101111010110111001001111111110111001100011111000101010";
                    when "01100" => level_vec_out <= "0101111100101111010110111001001111111111111001100011111000101010";
                    when "01101" => level_vec_out <= "0101111100101111010110111001001111111111111011100011111000101010";
                    when "01110" => level_vec_out <= "0101111100101111010110111001001111111111111011100111111000101010";
                    when "01111" => level_vec_out <= "0101111100101111010110111001001111111111111011100111111000101010";
                    when "10000" => level_vec_out <= "0101111100101111010110111001001111111111111011110111111000101010";
                    when "10001" => level_vec_out <= "0101111100101111110110111001001111111111111011111111111001101010";
                    when "10010" => level_vec_out <= "0101111100101111111110111001001111111111111011111111111001101010";
                    when "10011" => level_vec_out <= "0101111100101111111110111001001111111111111011111111111001101011";
                    when "10100" => level_vec_out <= "0101111100101111111110111011101111111111111011111111111001101011";
                    when "10101" => level_vec_out <= "0101111100101111111110111011101111111111111011111111111001101011";
                    when "10110" => level_vec_out <= "0101111100101111111110111111101111111111111011111111111011101011";
                    when "10111" => level_vec_out <= "0101111101101111111111111111101111111111111011111111111011101011";
                    when "11000" => level_vec_out <= "1101111101101111111111111111101111111111111011111111111011101011";
                    when "11001" => level_vec_out <= "1101111101101111111111111111101111111111111011111111111011101011";
                    when "11010" => level_vec_out <= "1111111101101111111111111111101111111111111011111111111011101011";
                    when "11011" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111011101011";
                    when "11100" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111011101011";
                    when "11101" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111011111011";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111011";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111011";
                when others => null;
                end case;
            when "101" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0111110000110100111011111100011110110011100100000110100111010110";
                    when "00001" => level_vec_out <= "0111110000110100111011111100011110110011100100000110100111010110";
                    when "00010" => level_vec_out <= "1111110000110100111011111100011110110011100100000110100111010110";
                    when "00011" => level_vec_out <= "1111110000111100111011111100011110110011100100000110100111010110";
                    when "00100" => level_vec_out <= "1111110000111100111011111101011110110011100100100110100111010110";
                    when "00101" => level_vec_out <= "1111110000111100111011111101011110110011100100110110100111010110";
                    when "00110" => level_vec_out <= "1111110000111101111011111101011110110011100100110110100111010110";
                    when "00111" => level_vec_out <= "1111110000111101111011111101111110110011100100110110100111010110";
                    when "01000" => level_vec_out <= "1111111000111101111011111101111110110011100100110110100111010110";
                    when "01001" => level_vec_out <= "1111111000111101111011111101111110110011100100111110100111010110";
                    when "01010" => level_vec_out <= "1111111000111101111011111101111110110011100100111110100111010110";
                    when "01011" => level_vec_out <= "1111111011111101111011111101111110110011100100111110100111010110";
                    when "01100" => level_vec_out <= "1111111011111101111011111101111110110011100101111110100111010110";
                    when "01101" => level_vec_out <= "1111111011111101111011111101111110110011100101111110110111010111";
                    when "01110" => level_vec_out <= "1111111011111101111011111101111110110011100101111110110111010111";
                    when "01111" => level_vec_out <= "1111111011111101111011111101111110110011101101111110110111010111";
                    when "10000" => level_vec_out <= "1111111011111101111111111101111110110111101101111110110111010111";
                    when "10001" => level_vec_out <= "1111111011111101111111111101111110111111101101111110110111010111";
                    when "10010" => level_vec_out <= "1111111011111101111111111101111110111111101101111110110111010111";
                    when "10011" => level_vec_out <= "1111111011111101111111111101111110111111101101111110110111110111";
                    when "10100" => level_vec_out <= "1111111011111101111111111101111110111111101101111111110111110111";
                    when "10101" => level_vec_out <= "1111111011111101111111111101111110111111111101111111110111110111";
                    when "10110" => level_vec_out <= "1111111011111101111111111101111110111111111101111111110111110111";
                    when "10111" => level_vec_out <= "1111111011111101111111111101111110111111111101111111110111110111";
                    when "11000" => level_vec_out <= "1111111011111101111111111101111110111111111101111111110111110111";
                    when "11001" => level_vec_out <= "1111111011111101111111111111111110111111111101111111110111110111";
                    when "11010" => level_vec_out <= "1111111011111101111111111111111110111111111101111111110111111111";
                    when "11011" => level_vec_out <= "1111111111111101111111111111111110111111111101111111110111111111";
                    when "11100" => level_vec_out <= "1111111111111101111111111111111110111111111101111111111111111111";
                    when "11101" => level_vec_out <= "1111111111111101111111111111111110111111111101111111111111111111";
                    when "11110" => level_vec_out <= "1111111111111101111111111111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "110" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1111100111011010001001101011010100110111100110101100100010101000";
                    when "00001" => level_vec_out <= "1111100111011010001001101011010100110111100110101100100010101100";
                    when "00010" => level_vec_out <= "1111100111011010001001101011010101110111100111101100100010101110";
                    when "00011" => level_vec_out <= "1111100111011010001001101011010101110111100111101101100010101110";
                    when "00100" => level_vec_out <= "1111100111011010001001101011110101110111100111101101100010101110";
                    when "00101" => level_vec_out <= "1111100111011010001001101011110101110111100111101101110110101110";
                    when "00110" => level_vec_out <= "1111100111011010001001101011110101110111100111101101110110101110";
                    when "00111" => level_vec_out <= "1111100111011010001001101011110111110111100111101101110110101110";
                    when "01000" => level_vec_out <= "1111100111011010001001101011110111110111110111111101110110101110";
                    when "01001" => level_vec_out <= "1111100111011010001001101011110111110111110111111101110110101110";
                    when "01010" => level_vec_out <= "1111100111011010001001101011110111110111110111111101110110101110";
                    when "01011" => level_vec_out <= "1111100111011010001001101011110111110111110111111111110110101110";
                    when "01100" => level_vec_out <= "1111100111111010001101111011110111110111110111111111110110101110";
                    when "01101" => level_vec_out <= "1111100111111010001101111011110111110111110111111111110110101110";
                    when "01110" => level_vec_out <= "1111100111111010001101111011110111110111110111111111110110101110";
                    when "01111" => level_vec_out <= "1111100111111010001101111011110111110111110111111111110110101110";
                    when "10000" => level_vec_out <= "1111100111111010001111111011110111110111110111111111110110101110";
                    when "10001" => level_vec_out <= "1111100111111010001111111011110111111111110111111111110110101110";
                    when "10010" => level_vec_out <= "1111100111111010001111111011110111111111110111111111110110101110";
                    when "10011" => level_vec_out <= "1111100111111010001111111011110111111111110111111111110110101110";
                    when "10100" => level_vec_out <= "1111100111111010001111111011110111111111111111111111110110111110";
                    when "10101" => level_vec_out <= "1111110111111010001111111011110111111111111111111111110110111110";
                    when "10110" => level_vec_out <= "1111110111111010001111111011110111111111111111111111110110111110";
                    when "10111" => level_vec_out <= "1111110111111010001111111011110111111111111111111111110110111110";
                    when "11000" => level_vec_out <= "1111110111111010001111111011110111111111111111111111110110111110";
                    when "11001" => level_vec_out <= "1111110111111010111111111011110111111111111111111111110111111110";
                    when "11010" => level_vec_out <= "1111110111111011111111111011110111111111111111111111110111111110";
                    when "11011" => level_vec_out <= "1111110111111011111111111011110111111111111111111111110111111110";
                    when "11100" => level_vec_out <= "1111110111111011111111111011110111111111111111111111111111111110";
                    when "11101" => level_vec_out <= "1111110111111011111111111111111111111111111111111111111111111110";
                    when "11110" => level_vec_out <= "1111110111111011111111111111111111111111111111111111111111111110";
                    when "11111" => level_vec_out <= "1111111111111011111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "111" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0110000010100110000110101100111000000011100000010101010001010101";
                    when "00001" => level_vec_out <= "0110000010100110010110101100111000000011100000010101010001010101";
                    when "00010" => level_vec_out <= "0110000010100110010110101100111000000011100000010101110001010101";
                    when "00011" => level_vec_out <= "0110000010100110010110101100111000000011100000010101110001010101";
                    when "00100" => level_vec_out <= "0110100010100110010110101100111000000011100000010101111001010101";
                    when "00101" => level_vec_out <= "0110100010100110010110101100111000000011100000010101111001010101";
                    when "00110" => level_vec_out <= "0110100010100110010110101100111000000011100000010101111001010101";
                    when "00111" => level_vec_out <= "0110100010100110010110101100111000000011100000010101111001010101";
                    when "01000" => level_vec_out <= "0110110010100110010110101100111000000011100000010101111001010101";
                    when "01001" => level_vec_out <= "0110110010100110010110101100111010000011100000010101111001010101";
                    when "01010" => level_vec_out <= "0110110010101110010110101100111010000011100000110101111001010101";
                    when "01011" => level_vec_out <= "0110110010101110110110101100111010010011100010110101111001010101";
                    when "01100" => level_vec_out <= "0110110010101111110110101100111010010011100110110101111001010101";
                    when "01101" => level_vec_out <= "0110110010101111110110101100111010010011100110110101111001010101";
                    when "01110" => level_vec_out <= "0110110010101111110110101101111010010011100110110101111001010101";
                    when "01111" => level_vec_out <= "0111110010101111110111101101111010010011100110110101111001010101";
                    when "10000" => level_vec_out <= "0111110010101111110111101101111010010011100110110101111001011101";
                    when "10001" => level_vec_out <= "0111110010101111110111101101111010010011100110110101111001011101";
                    when "10010" => level_vec_out <= "0111110010101111110111111111111010010011100110110101111001011101";
                    when "10011" => level_vec_out <= "0111110010101111110111111111111010110011100110110101111001011101";
                    when "10100" => level_vec_out <= "0111111010101111110111111111111010110011100110110101111001011101";
                    when "10101" => level_vec_out <= "0111111010101111110111111111111010111011100110110101111011011101";
                    when "10110" => level_vec_out <= "0111111010101111110111111111111110111011100110110101111011011101";
                    when "10111" => level_vec_out <= "0111111010111111110111111111111110111011101110110101111011111101";
                    when "11000" => level_vec_out <= "0111111110111111110111111111111110111111101110110111111011111111";
                    when "11001" => level_vec_out <= "0111111110111111111111111111111110111111101110110111111011111111";
                    when "11010" => level_vec_out <= "0111111110111111111111111111111110111111111110110111111011111111";
                    when "11011" => level_vec_out <= "1111111111111111111111111111111110111111111110110111111011111111";
                    when "11100" => level_vec_out <= "1111111111111111111111111111111110111111111111111111111011111111";
                    when "11101" => level_vec_out <= "1111111111111111111111111111111110111111111111111111111011111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111110111111111111111111111011111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when others => null;
        end case;
    end process;
end Behavioral;