----
 -- @file level_hvec_gen_hdl.hpp
 -- @brief This script generates HDL code for generating high-dimensional LEVEL vectors.
 -- It is a novel method; for more information, please refer to our paper.
 --
 -- @author Saeid Jamili and Marco Angioli
 -- @note Author names are listed in alphabetical order.
 -- @email <saeid.jamili@uniroma1.it>
 -- @email <marco.angioli@uniroma1.it>
 --
 -- @contributors
 --
 -- @date Created: 24th July 2023
 -- @date Last Updated: 23th August 2023
 --
 -- @version 1.0.0
 --
 -- @institute Sapienza University of Rome
 -- @cite https://doi.org/10.xxxx/yyyyy
 --
 -- @section DEPENDENCIES
 -- - Dependency1: Description or version details.
 -- - Dependency2: Description or version details.
 --
 -- @section LICENSE
 -- This file is part of the Aeneas HyperCompute Platform.
 --
 -- Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 --
 -- @section CHANGELOG
 -- @version 1.0.0-dev - 23th August 2023
 -- - Initial release
 --
 -- @todo
 -- - Complete level vector generator function
 -- - Add training
 --
 -- @see
 -- -
 -- -
 -- -
 --
 --

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity level_vec_gen is
    Port ( level_vec_out : out  STD_LOGIC_VECTOR (63 downto 0);
           frame_index : in  STD_LOGIC_VECTOR (2 downto 0);
           frame_id : in  STD_LOGIC_VECTOR (4 downto 0));
end level_vec_gen;

architecture Behavioral of level_vec_gen is
begin
    process (frame_index, frame_id)
    begin
        -- Update this function to match your requirements
        case frame_index is
            when "000" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00001" => level_vec_out <= "1111111111111111000000000000000000000000000000000000000000000000";
                    when "00010" => level_vec_out <= "1111111111111111111111110000000000000000000000000000000000000000";
                    when "00011" => level_vec_out <= "1111111111111111111111111111111100000000000000000000000000000000";
                    when "00100" => level_vec_out <= "1111111111111111111111111111111111111111000000000000000000000000";
                    when "00101" => level_vec_out <= "1111111111111111111111111111111111111111111111110000000000000000";
                    when "00110" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111100000000";
                    when "00111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "01000" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "01001" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "01010" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "01011" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "01100" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "01101" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "01110" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "01111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "10000" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "10001" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "10010" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "10011" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "10100" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "10101" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "10110" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "10111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "11000" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "11001" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "11010" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "11011" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "11100" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "11101" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "001" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00001" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00010" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00011" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00100" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00101" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00110" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00111" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "01000" => level_vec_out <= "1111111100000000000000000000000000000000000000000000000000000000";
                    when "01001" => level_vec_out <= "1111111111111111000000000000000000000000000000000000000000000000";
                    when "01010" => level_vec_out <= "1111111111111111111111110000000000000000000000000000000000000000";
                    when "01011" => level_vec_out <= "1111111111111111111111111111111100000000000000000000000000000000";
                    when "01100" => level_vec_out <= "1111111111111111111111111111111111111111000000000000000000000000";
                    when "01101" => level_vec_out <= "1111111111111111111111111111111111111111111111110000000000000000";
                    when "01110" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111100000000";
                    when "01111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "10000" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "10001" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "10010" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "10011" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "10100" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "10101" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "10110" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "10111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "11000" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "11001" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "11010" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "11011" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "11100" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "11101" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "010" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00001" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00010" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00011" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00100" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00101" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00110" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00111" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "01000" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "01001" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "01010" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "01011" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "01100" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "01101" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "01110" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "01111" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "10000" => level_vec_out <= "1111111100000000000000000000000000000000000000000000000000000000";
                    when "10001" => level_vec_out <= "1111111111111111000000000000000000000000000000000000000000000000";
                    when "10010" => level_vec_out <= "1111111111111111111111110000000000000000000000000000000000000000";
                    when "10011" => level_vec_out <= "1111111111111111111111111111111100000000000000000000000000000000";
                    when "10100" => level_vec_out <= "1111111111111111111111111111111111111111000000000000000000000000";
                    when "10101" => level_vec_out <= "1111111111111111111111111111111111111111111111110000000000000000";
                    when "10110" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111100000000";
                    when "10111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "11000" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "11001" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "11010" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "11011" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "11100" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "11101" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "011" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00001" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00010" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00011" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00100" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00101" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00110" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00111" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "01000" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "01001" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "01010" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "01011" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "01100" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "01101" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "01110" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "01111" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "10000" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "10001" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "10010" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "10011" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "10100" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "10101" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "10110" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "10111" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "11000" => level_vec_out <= "1111111100000000000000000000000000000000000000000000000000000000";
                    when "11001" => level_vec_out <= "1111111111111111000000000000000000000000000000000000000000000000";
                    when "11010" => level_vec_out <= "1111111111111111111111110000000000000000000000000000000000000000";
                    when "11011" => level_vec_out <= "1111111111111111111111111111111100000000000000000000000000000000";
                    when "11100" => level_vec_out <= "1111111111111111111111111111111111111111000000000000000000000000";
                    when "11101" => level_vec_out <= "1111111111111111111111111111111111111111111111110000000000000000";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111100000000";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "100" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00001" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00010" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00011" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00100" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00101" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00110" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00111" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "01000" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "01001" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "01010" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "01011" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "01100" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "01101" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "01110" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "01111" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "10000" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "10001" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "10010" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "10011" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "10100" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "10101" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "10110" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "10111" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "11000" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "11001" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "11010" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "11011" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "11100" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "11101" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "11110" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "11111" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                when others => null;
                end case;
            when "101" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00001" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00010" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00011" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00100" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00101" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00110" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00111" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "01000" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "01001" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "01010" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "01011" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "01100" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "01101" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "01110" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "01111" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "10000" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "10001" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "10010" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "10011" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "10100" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "10101" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "10110" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "10111" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "11000" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "11001" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "11010" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "11011" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "11100" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "11101" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "11110" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "11111" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                when others => null;
                end case;
            when "110" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00001" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00010" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00011" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00100" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00101" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00110" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00111" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "01000" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "01001" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "01010" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "01011" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "01100" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "01101" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "01110" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "01111" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "10000" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "10001" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "10010" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "10011" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "10100" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "10101" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "10110" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "10111" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "11000" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "11001" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "11010" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "11011" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "11100" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "11101" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "11110" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "11111" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                when others => null;
                end case;
            when "111" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00001" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00010" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00011" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00100" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00101" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00110" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "00111" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "01000" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "01001" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "01010" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "01011" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "01100" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "01101" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "01110" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "01111" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "10000" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "10001" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "10010" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "10011" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "10100" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "10101" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "10110" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "10111" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "11000" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "11001" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "11010" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "11011" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "11100" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "11101" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "11110" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                    when "11111" => level_vec_out <= "0000000000000000000000000000000000000000000000000000000000000000";
                when others => null;
                end case;
            when others => null;
        end case;
    end process;
end Behavioral;