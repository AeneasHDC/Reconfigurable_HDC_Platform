/**
 * @file level_hvec_gen_hdl.hpp
 * @brief This script generates HDL code for generating high-dimensional LEVEL vectors.
 * It is a novel method; for more information, please refer to our paper.
 *
 * @author Saeid Jamili and Marco Angioli
 * @note Author names are listed in alphabetical order.
 * @email <saeid.jamili@uniroma1.it>
 * @email <marco.angioli@uniroma1.it>
 *
 * @contributors
 *
 * @date Created: 24th July 2023
 * @date Last Updated: 23th August 2023
 *
 * @version 1.0.0
 *
 * @institute Sapienza University of Rome
 * @cite https://doi.org/10.xxxx/yyyyy
 *
 * @section DEPENDENCIES
 * - Dependency1: Description or version details.
 * - Dependency2: Description or version details.
 *
 * @section LICENSE
 * This file is part of the Aeneas HyperCompute Platform.
 *
 * Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 *
 * @section CHANGELOG
 * @version 1.0.0-dev - 23th August 2023
 * - Initial release
 *
 * @todo
 * - Complete level vector generator function
 * - Add training
 *
 * @see
 * -
 * -
 * -
 *
 */

module level_vec_gen (
    output reg [63:0] level_vec_out,
    input [2:0] frame_index,
    input [4:0] frame_id
);
    always @(*) begin
        // Update this function to match your requirements
        case (frame_index)
            0: begin
                case (frame_id)
                    0: level_vec_out = 64'b1110000000001001111110100000001000001011111110001010101010101100;
                    1: level_vec_out = 64'b1110000000001001111110100000001000001011111111001010101010101100;
                    2: level_vec_out = 64'b1110000000001001111110100000001000001011111111001010101010101100;
                    3: level_vec_out = 64'b1110000000001001111110100000001010001011111111001010111010101100;
                    4: level_vec_out = 64'b1110000000001001111110100000001010001011111111101010111010101100;
                    5: level_vec_out = 64'b1110000000001001111110100000001010001011111111101010111010101100;
                    6: level_vec_out = 64'b1110000100001001111110100000001010001011111111111010111010101100;
                    7: level_vec_out = 64'b1110000100001001111110100000001010001011111111111010111010101100;
                    8: level_vec_out = 64'b1111000100001001111110100000001010001011111111111110111010101100;
                    9: level_vec_out = 64'b1111000100001101111110100000001010001011111111111110111010101100;
                    10: level_vec_out = 64'b1111000100001101111110100000001010001011111111111110111010111100;
                    11: level_vec_out = 64'b1111000100101101111110100000001010001011111111111110111010111101;
                    12: level_vec_out = 64'b1111000100101101111111110000001010001011111111111110111010111101;
                    13: level_vec_out = 64'b1111000100101101111111110000001010001011111111111111111010111101;
                    14: level_vec_out = 64'b1111000100101101111111110000001010001011111111111111111010111101;
                    15: level_vec_out = 64'b1111000100101101111111110000001010001011111111111111111010111101;
                    16: level_vec_out = 64'b1111100100101101111111111000001010001011111111111111111110111101;
                    17: level_vec_out = 64'b1111100100101101111111111000001010101011111111111111111110111101;
                    18: level_vec_out = 64'b1111100100101101111111111000011010101011111111111111111110111111;
                    19: level_vec_out = 64'b1111101100101111111111111000011010101111111111111111111110111111;
                    20: level_vec_out = 64'b1111101100101111111111111001011010101111111111111111111110111111;
                    21: level_vec_out = 64'b1111101100101111111111111001111010101111111111111111111111111111;
                    22: level_vec_out = 64'b1111101100101111111111111001111011101111111111111111111111111111;
                    23: level_vec_out = 64'b1111101100101111111111111101111011101111111111111111111111111111;
                    24: level_vec_out = 64'b1111101100101111111111111101111011101111111111111111111111111111;
                    25: level_vec_out = 64'b1111101100101111111111111101111111101111111111111111111111111111;
                    26: level_vec_out = 64'b1111111100101111111111111111111111101111111111111111111111111111;
                    27: level_vec_out = 64'b1111111100101111111111111111111111101111111111111111111111111111;
                    28: level_vec_out = 64'b1111111100101111111111111111111111101111111111111111111111111111;
                    29: level_vec_out = 64'b1111111100101111111111111111111111101111111111111111111111111111;
                    30: level_vec_out = 64'b1111111110111111111111111111111111111111111111111111111111111111;
                    31: level_vec_out = 64'b1111111110111111111111111111111111111111111111111111111111111111;
                endcase
            end
            1: begin
                case (frame_id)
                    0: level_vec_out = 64'b1001111011001110000101100000010000101110100001010101011010000001;
                    1: level_vec_out = 64'b1001111011001110000101100000010000101110100001010101011010000001;
                    2: level_vec_out = 64'b1001111011001110001101100000010000101110100001010101011011000001;
                    3: level_vec_out = 64'b1001111011001110001101100000010000101110100001010101111011000001;
                    4: level_vec_out = 64'b1001111011001110001101100000010000101110100001010101111011000001;
                    5: level_vec_out = 64'b1001111011001110001101100000010000101110100001010101111011000001;
                    6: level_vec_out = 64'b1001111011001110001101100010010000101110100001011101111011100001;
                    7: level_vec_out = 64'b1101111011001110001101100010010010101110100001011101111011100001;
                    8: level_vec_out = 64'b1101111011001110001101100010010010101110100001011101111011100001;
                    9: level_vec_out = 64'b1101111011001110101101100110010010101110100001011101111011100001;
                    10: level_vec_out = 64'b1101111011001110101111100110010010101110100001011101111011100001;
                    11: level_vec_out = 64'b1101111011001110101111100111010010101110100001011101111011100001;
                    12: level_vec_out = 64'b1101111011001110101111110111011010101110100001011101111011100001;
                    13: level_vec_out = 64'b1101111011001110101111110111011010101110100011011101111011100001;
                    14: level_vec_out = 64'b1101111011001110101111110111111010101110100011011101111011100001;
                    15: level_vec_out = 64'b1101111011001110111111110111111010101110110011011101111011100001;
                    16: level_vec_out = 64'b1101111011001110111111110111111010101110110011111101111011100001;
                    17: level_vec_out = 64'b1101111011001110111111110111111010101110111011111101111011100001;
                    18: level_vec_out = 64'b1101111011011110111111110111111010101110111011111101111111100001;
                    19: level_vec_out = 64'b1101111011011110111111110111111010111110111011111101111111100001;
                    20: level_vec_out = 64'b1101111011011110111111110111111010111110111011111101111111100001;
                    21: level_vec_out = 64'b1101111011011110111111110111111010111110111111111101111111100001;
                    22: level_vec_out = 64'b1101111011011110111111111111111010111110111111111101111111100101;
                    23: level_vec_out = 64'b1111111011011110111111111111111011111110111111111101111111100101;
                    24: level_vec_out = 64'b1111111011011110111111111111111011111111111111111101111111100101;
                    25: level_vec_out = 64'b1111111011011111111111111111111011111111111111111101111111100111;
                    26: level_vec_out = 64'b1111111011011111111111111111111011111111111111111101111111110111;
                    27: level_vec_out = 64'b1111111111011111111111111111111011111111111111111101111111110111;
                    28: level_vec_out = 64'b1111111111111111111111111111111111111111111111111101111111110111;
                    29: level_vec_out = 64'b1111111111111111111111111111111111111111111111111101111111110111;
                    30: level_vec_out = 64'b1111111111111111111111111111111111111111111111111101111111110111;
                    31: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111110111;
                endcase
            end
            2: begin
                case (frame_id)
                    0: level_vec_out = 64'b1010011000011111110011011111100011001010110111101011001011000000;
                    1: level_vec_out = 64'b1010011000011111110011011111100011001010110111101011001011000000;
                    2: level_vec_out = 64'b1010011000011111110011011111100011001010111111101011001011000000;
                    3: level_vec_out = 64'b1010011000011111110011011111100011001010111111101011001011000000;
                    4: level_vec_out = 64'b1010011000011111110011011111100011001010111111101011001011000000;
                    5: level_vec_out = 64'b1010011000011111110011011111100011001010111111101011001111000000;
                    6: level_vec_out = 64'b1010011000011111110011011111100011001010111111111011001111001000;
                    7: level_vec_out = 64'b1010011000011111110011011111100011001010111111111011001111001010;
                    8: level_vec_out = 64'b1011011000011111110011111111100011001010111111111111001111001010;
                    9: level_vec_out = 64'b1011011000011111110011111111100011001010111111111111001111001010;
                    10: level_vec_out = 64'b1011011000011111110011111111100011001010111111111111001111001010;
                    11: level_vec_out = 64'b1011011000011111111011111111100011001010111111111111001111001010;
                    12: level_vec_out = 64'b1011111000011111111011111111100011001110111111111111001111001010;
                    13: level_vec_out = 64'b1011111000011111111011111111100011001110111111111111001111001010;
                    14: level_vec_out = 64'b1011111000011111111011111111100011011110111111111111001111001010;
                    15: level_vec_out = 64'b1011111000111111111111111111100011011110111111111111001111001010;
                    16: level_vec_out = 64'b1011111100111111111111111111100011011110111111111111001111001010;
                    17: level_vec_out = 64'b1011111100111111111111111111100011011110111111111111001111001010;
                    18: level_vec_out = 64'b1011111100111111111111111111100011011110111111111111001111001010;
                    19: level_vec_out = 64'b1011111101111111111111111111100111011110111111111111001111001010;
                    20: level_vec_out = 64'b1011111101111111111111111111110111011110111111111111011111001010;
                    21: level_vec_out = 64'b1111111111111111111111111111110111011110111111111111011111001010;
                    22: level_vec_out = 64'b1111111111111111111111111111110111111110111111111111011111101010;
                    23: level_vec_out = 64'b1111111111111111111111111111110111111110111111111111011111101110;
                    24: level_vec_out = 64'b1111111111111111111111111111111111111110111111111111011111101110;
                    25: level_vec_out = 64'b1111111111111111111111111111111111111110111111111111011111101110;
                    26: level_vec_out = 64'b1111111111111111111111111111111111111110111111111111011111101110;
                    27: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111011111111110;
                    28: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111110;
                    29: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111110;
                    30: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111110;
                    31: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111110;
                endcase
            end
            3: begin
                case (frame_id)
                    0: level_vec_out = 64'b0011010011100110000001011101111111100011011011100001110111111000;
                    1: level_vec_out = 64'b0011010011100110000001011101111111100011011111100001110111111000;
                    2: level_vec_out = 64'b0011010011100110001001011101111111100011011111100001110111111000;
                    3: level_vec_out = 64'b0011010011101110001001011101111111100011011111100001110111111000;
                    4: level_vec_out = 64'b0011010011101110001001011101111111100011011111100001110111111000;
                    5: level_vec_out = 64'b0011010011101110001001011101111111110011011111100011110111111000;
                    6: level_vec_out = 64'b0011010011101110001001011101111111110011011111100011110111111000;
                    7: level_vec_out = 64'b0011010011101110001001011101111111110111011111100011110111111000;
                    8: level_vec_out = 64'b0011010011101110001001011101111111110111011111100011110111111000;
                    9: level_vec_out = 64'b0011010011101110001001011101111111111111011111100011110111111000;
                    10: level_vec_out = 64'b0011010011101110001001011101111111111111011111100011110111111001;
                    11: level_vec_out = 64'b0011011011101110001001011101111111111111011111100011110111111001;
                    12: level_vec_out = 64'b0011011011101110001001011101111111111111011111100011110111111011;
                    13: level_vec_out = 64'b0011011011101110001001011101111111111111011111100011110111111011;
                    14: level_vec_out = 64'b0011011011101110011001011101111111111111011111100011110111111011;
                    15: level_vec_out = 64'b0011011011101111011001011101111111111111011111100011110111111011;
                    16: level_vec_out = 64'b0011111011101111011001011101111111111111011111100011110111111011;
                    17: level_vec_out = 64'b0011111011101111011001011101111111111111111111101011110111111011;
                    18: level_vec_out = 64'b0011111011101111011001011111111111111111111111101011110111111011;
                    19: level_vec_out = 64'b0011111011101111011001011111111111111111111111101011110111111011;
                    20: level_vec_out = 64'b0111111011101111011001011111111111111111111111101011110111111011;
                    21: level_vec_out = 64'b0111111011101111011001011111111111111111111111101011110111111011;
                    22: level_vec_out = 64'b0111111011101111011001011111111111111111111111101011110111111011;
                    23: level_vec_out = 64'b0111111011101111011001011111111111111111111111101011110111111011;
                    24: level_vec_out = 64'b0111111011101111011001011111111111111111111111101011110111111011;
                    25: level_vec_out = 64'b0111111011101111011001011111111111111111111111101011110111111011;
                    26: level_vec_out = 64'b0111111011101111011101011111111111111111111111101011110111111011;
                    27: level_vec_out = 64'b0111111011101111011111011111111111111111111111101011110111111111;
                    28: level_vec_out = 64'b0111111011111111011111011111111111111111111111101011110111111111;
                    29: level_vec_out = 64'b1111111011111111011111111111111111111111111111101011111111111111;
                    30: level_vec_out = 64'b1111111111111111011111111111111111111111111111101111111111111111;
                    31: level_vec_out = 64'b1111111111111111111111111111111111111111111111101111111111111111;
                endcase
            end
            4: begin
                case (frame_id)
                    0: level_vec_out = 64'b1100010101100100110101010000010101000111111110100011100001011110;
                    1: level_vec_out = 64'b1100010101100100110101110000010101000111111110100011100001011110;
                    2: level_vec_out = 64'b1110010101100100110101110000010101000111111111100011100001011110;
                    3: level_vec_out = 64'b1110010101100110110101110000010101000111111111100011100001011110;
                    4: level_vec_out = 64'b1110010101101110110101110000010111000111111111100111100001011110;
                    5: level_vec_out = 64'b1110010101101110110101110000010111000111111111100111100001011110;
                    6: level_vec_out = 64'b1110010101101110110101110000010111000111111111100111100001011110;
                    7: level_vec_out = 64'b1110010101101110110101110000010111000111111111100111101001011110;
                    8: level_vec_out = 64'b1110010101101110110101110000110111000111111111100111101001011110;
                    9: level_vec_out = 64'b1110010101101110110101110001110111000111111111100111101001011110;
                    10: level_vec_out = 64'b1110010101101110110101110001110111010111111111100111101001011110;
                    11: level_vec_out = 64'b1110010101101110110101110001110111010111111111100111101001011110;
                    12: level_vec_out = 64'b1110010101101110110101110001110111010111111111100111101001011110;
                    13: level_vec_out = 64'b1110010101101110110101110001110111010111111111100111101001011110;
                    14: level_vec_out = 64'b1110010101101110110101110001110111010111111111100111101001011111;
                    15: level_vec_out = 64'b1110010101101110110111110001110111010111111111101111101001011111;
                    16: level_vec_out = 64'b1110110101101110110111110001110111010111111111101111101001011111;
                    17: level_vec_out = 64'b1110110101101111110111110001110111010111111111101111101001111111;
                    18: level_vec_out = 64'b1110110101101111110111110001110111010111111111101111101001111111;
                    19: level_vec_out = 64'b1110110101101111110111110001110111010111111111101111101001111111;
                    20: level_vec_out = 64'b1110110101101111110111110001110111010111111111101111111001111111;
                    21: level_vec_out = 64'b1110110111101111110111110001110111010111111111101111111001111111;
                    22: level_vec_out = 64'b1110110111101111110111110001110111110111111111101111111001111111;
                    23: level_vec_out = 64'b1111110111101111110111110001110111110111111111101111111001111111;
                    24: level_vec_out = 64'b1111110111101111110111110001110111110111111111111111111001111111;
                    25: level_vec_out = 64'b1111110111101111110111111001110111110111111111111111111001111111;
                    26: level_vec_out = 64'b1111110111101111111111111001110111110111111111111111111001111111;
                    27: level_vec_out = 64'b1111110111101111111111111001110111110111111111111111111001111111;
                    28: level_vec_out = 64'b1111111111101111111111111101110111110111111111111111111001111111;
                    29: level_vec_out = 64'b1111111111111111111111111101111111110111111111111111111101111111;
                    30: level_vec_out = 64'b1111111111111111111111111101111111110111111111111111111101111111;
                    31: level_vec_out = 64'b1111111111111111111111111111111111110111111111111111111101111111;
                endcase
            end
            5: begin
                case (frame_id)
                    0: level_vec_out = 64'b1011001100000001101101111111100010010101000101100110101111010111;
                    1: level_vec_out = 64'b1111001100000001101101111111111010010101000101100110101111010111;
                    2: level_vec_out = 64'b1111001100000001101101111111111010010101000101100110101111010111;
                    3: level_vec_out = 64'b1111001100000001101101111111111010010101001101100110101111010111;
                    4: level_vec_out = 64'b1111001110000001101101111111111010010101001101100110101111010111;
                    5: level_vec_out = 64'b1111001110010001101101111111111010010101001101100111101111010111;
                    6: level_vec_out = 64'b1111001110010001101101111111111010010101001101100111111111010111;
                    7: level_vec_out = 64'b1111001111110001101101111111111010010101001101100111111111010111;
                    8: level_vec_out = 64'b1111001111110001101101111111111010010101001101100111111111010111;
                    9: level_vec_out = 64'b1111001111110001111101111111111010010101001101100111111111010111;
                    10: level_vec_out = 64'b1111001111110001111101111111111010010101001101100111111111110111;
                    11: level_vec_out = 64'b1111101111110001111101111111111010010101001101100111111111110111;
                    12: level_vec_out = 64'b1111101111110001111101111111111010010101101101100111111111110111;
                    13: level_vec_out = 64'b1111101111110001111101111111111010010101101101100111111111110111;
                    14: level_vec_out = 64'b1111101111110001111101111111111110010101101101101111111111111111;
                    15: level_vec_out = 64'b1111101111110001111101111111111110010101101101101111111111111111;
                    16: level_vec_out = 64'b1111101111110001111101111111111110010101101101101111111111111111;
                    17: level_vec_out = 64'b1111101111110001111101111111111110010101101101101111111111111111;
                    18: level_vec_out = 64'b1111101111110001111101111111111110010101101101111111111111111111;
                    19: level_vec_out = 64'b1111101111110001111101111111111110010101101101111111111111111111;
                    20: level_vec_out = 64'b1111101111110101111101111111111110010111101101111111111111111111;
                    21: level_vec_out = 64'b1111101111110101111101111111111111010111101101111111111111111111;
                    22: level_vec_out = 64'b1111101111110101111101111111111111010111101101111111111111111111;
                    23: level_vec_out = 64'b1111101111110101111101111111111111010111101101111111111111111111;
                    24: level_vec_out = 64'b1111101111111101111101111111111111010111101101111111111111111111;
                    25: level_vec_out = 64'b1111101111111101111101111111111111111111101101111111111111111111;
                    26: level_vec_out = 64'b1111101111111101111101111111111111111111111111111111111111111111;
                    27: level_vec_out = 64'b1111101111111101111111111111111111111111111111111111111111111111;
                    28: level_vec_out = 64'b1111101111111111111111111111111111111111111111111111111111111111;
                    29: level_vec_out = 64'b1111101111111111111111111111111111111111111111111111111111111111;
                    30: level_vec_out = 64'b1111101111111111111111111111111111111111111111111111111111111111;
                    31: level_vec_out = 64'b1111101111111111111111111111111111111111111111111111111111111111;
                endcase
            end
            6: begin
                case (frame_id)
                    0: level_vec_out = 64'b0001111111111000111001111111011101110100110010101001100010001110;
                    1: level_vec_out = 64'b0001111111111000111001111111111101110101110010101001100010001110;
                    2: level_vec_out = 64'b0001111111111000111001111111111101110101110010101001100010001110;
                    3: level_vec_out = 64'b0001111111111000111001111111111101110101110010101001100010011111;
                    4: level_vec_out = 64'b0001111111111010111001111111111101110101110010101011100010011111;
                    5: level_vec_out = 64'b0001111111111010111001111111111101110101110011101011100010011111;
                    6: level_vec_out = 64'b0001111111111010111001111111111101110101110011101011100010011111;
                    7: level_vec_out = 64'b0001111111111010111001111111111101110101110011101011100010011111;
                    8: level_vec_out = 64'b0001111111111110111001111111111101110101110111101011100010011111;
                    9: level_vec_out = 64'b0001111111111110111101111111111101110101110111101011100010011111;
                    10: level_vec_out = 64'b0001111111111111111101111111111111110101110111101011100010011111;
                    11: level_vec_out = 64'b0001111111111111111101111111111111110111110111101011100010011111;
                    12: level_vec_out = 64'b0001111111111111111101111111111111110111110111101011100010011111;
                    13: level_vec_out = 64'b0101111111111111111101111111111111111111111111101011100010011111;
                    14: level_vec_out = 64'b0101111111111111111101111111111111111111111111101011100010011111;
                    15: level_vec_out = 64'b0101111111111111111101111111111111111111111111101011100110011111;
                    16: level_vec_out = 64'b0101111111111111111101111111111111111111111111101011100110011111;
                    17: level_vec_out = 64'b0101111111111111111101111111111111111111111111101011100110011111;
                    18: level_vec_out = 64'b0101111111111111111101111111111111111111111111101111100110011111;
                    19: level_vec_out = 64'b0101111111111111111101111111111111111111111111101111110110011111;
                    20: level_vec_out = 64'b0101111111111111111101111111111111111111111111101111110110011111;
                    21: level_vec_out = 64'b0101111111111111111101111111111111111111111111101111111110011111;
                    22: level_vec_out = 64'b0101111111111111111101111111111111111111111111101111111111111111;
                    23: level_vec_out = 64'b1111111111111111111101111111111111111111111111101111111111111111;
                    24: level_vec_out = 64'b1111111111111111111101111111111111111111111111101111111111111111;
                    25: level_vec_out = 64'b1111111111111111111101111111111111111111111111101111111111111111;
                    26: level_vec_out = 64'b1111111111111111111101111111111111111111111111101111111111111111;
                    27: level_vec_out = 64'b1111111111111111111101111111111111111111111111101111111111111111;
                    28: level_vec_out = 64'b1111111111111111111101111111111111111111111111101111111111111111;
                    29: level_vec_out = 64'b1111111111111111111101111111111111111111111111101111111111111111;
                    30: level_vec_out = 64'b1111111111111111111101111111111111111111111111101111111111111111;
                    31: level_vec_out = 64'b1111111111111111111101111111111111111111111111111111111111111111;
                endcase
            end
            7: begin
                case (frame_id)
                    0: level_vec_out = 64'b0000101101001010001100110110000000000110011000000011100111101010;
                    1: level_vec_out = 64'b0000101101001010001100110110000000000110011000000011100111101010;
                    2: level_vec_out = 64'b0000101101001010001100110110000010000110011000000111100111101010;
                    3: level_vec_out = 64'b0000101101001010001100110110000010000110011000000111100111101010;
                    4: level_vec_out = 64'b0000101101001010001100110110010010000110011000000111100111101010;
                    5: level_vec_out = 64'b0000111101001010001100110110010010000110111000000111100111101010;
                    6: level_vec_out = 64'b0000111101001010001100110110010010000110111000000111100111101010;
                    7: level_vec_out = 64'b0000111101011010001100110110010010000110111000000111100111101010;
                    8: level_vec_out = 64'b0000111101011010001100110110010010000110111000000111100111101010;
                    9: level_vec_out = 64'b0000111101011010001100110110010010000110111000000111100111101110;
                    10: level_vec_out = 64'b0000111101011010001100110110010010000111111000000111100111101110;
                    11: level_vec_out = 64'b0000111101011010001100110110010010010111111000000111100111101110;
                    12: level_vec_out = 64'b0000111101011010001100110110010010010111111000000111100111101110;
                    13: level_vec_out = 64'b1000111101011010001100110110011010010111111000000111101111101110;
                    14: level_vec_out = 64'b1000111101011010001100110110011010010111111000010111101111101110;
                    15: level_vec_out = 64'b1000111101011010001100110110011010010111111000010111101111101110;
                    16: level_vec_out = 64'b1000111101011010001100111110011010010111111000010111101111101110;
                    17: level_vec_out = 64'b1000111101011010001110111110111010010111111000010111101111101110;
                    18: level_vec_out = 64'b1000111101011010001110111110111010010111111000010111101111111110;
                    19: level_vec_out = 64'b1000111101011010001110111110111010110111111000010111101111111110;
                    20: level_vec_out = 64'b1000111101011010001110111110111010110111111001010111101111111110;
                    21: level_vec_out = 64'b1000111101011010001110111110111010110111111001010111101111111110;
                    22: level_vec_out = 64'b1000111101011010001110111110111010110111111001010111101111111110;
                    23: level_vec_out = 64'b1000111101011010101110111110111010110111111001010111101111111110;
                    24: level_vec_out = 64'b1010111111111010111110111110111010110111111001010111101111111110;
                    25: level_vec_out = 64'b1011111111111010111110111111111010110111111001010111101111111110;
                    26: level_vec_out = 64'b1111111111111010111110111111111010110111111001010111101111111110;
                    27: level_vec_out = 64'b1111111111111111111110111111111010110111111001010111101111111110;
                    28: level_vec_out = 64'b1111111111111111111110111111111010110111111001010111101111111111;
                    29: level_vec_out = 64'b1111111111111111111110111111111010110111111001011111111111111111;
                    30: level_vec_out = 64'b1111111111111111111111111111111011110111111101011111111111111111;
                    31: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                endcase
            end
        endcase
    end
endmodule