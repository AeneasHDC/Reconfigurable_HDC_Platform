----
 -- @file level_hvec_gen_hdl.hpp
 -- @brief This script generates HDL code for generating high-dimensional LEVEL vectors.
 -- It is a novel method; for more information, please refer to our paper.
 --
 -- @author Saeid Jamili and Marco Angioli
 -- @note Author names are listed in alphabetical order.
 -- @email <saeid.jamili@uniroma1.it>
 -- @email <marco.angioli@uniroma1.it>
 --
 -- @contributors
 --
 -- @date Created: 24th July 2023
 -- @date Last Updated: 23th August 2023
 --
 -- @version 1.0.0
 --
 -- @institute Sapienza University of Rome
 -- @cite https://doi.org/10.xxxx/yyyyy
 --
 -- @section DEPENDENCIES
 -- - Dependency1: Description or version details.
 -- - Dependency2: Description or version details.
 --
 -- @section LICENSE
 -- This file is part of the Aeneas HyperCompute Platform.
 --
 -- Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 --
 -- @section CHANGELOG
 -- @version 1.0.0-dev - 23th August 2023
 -- - Initial release
 --
 -- @todo
 -- - Complete level vector generator function
 -- - Add training
 --
 -- @see
 -- -
 -- -
 -- -
 --
 --

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity level_vec_gen is
    Port ( level_vec_out : out  STD_LOGIC_VECTOR (63 downto 0);
           frame_index : in  STD_LOGIC_VECTOR (2 downto 0);
           frame_id : in  STD_LOGIC_VECTOR (4 downto 0));
end level_vec_gen;

architecture Behavioral of level_vec_gen is
begin
    process (frame_index, frame_id)
    begin
        -- Update this function to match your requirements
        case frame_index is
            when "000" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0000110101011001011101011011100100010001111010101101000100100000";
                    when "00001" => level_vec_out <= "1000110101011001011101111011100100010001111010101101000100100000";
                    when "00010" => level_vec_out <= "1000111101011001011101111011100100010001111010111101000100100000";
                    when "00011" => level_vec_out <= "1000111101011001011101111011100100010001111010111101000100100010";
                    when "00100" => level_vec_out <= "1000111101011011011111111011100100010001111010111101000100100010";
                    when "00101" => level_vec_out <= "1000111101011011011111111011110100010001111010111101000100100010";
                    when "00110" => level_vec_out <= "1000111101011011011111111011110100010001111110111111000100100010";
                    when "00111" => level_vec_out <= "1000111101011011011111111011110101011001111110111111000100100010";
                    when "01000" => level_vec_out <= "1000111101011011011111111011110101011001111110111111000100100010";
                    when "01001" => level_vec_out <= "1000111101011011011111111011110101011001111110111111000100100010";
                    when "01010" => level_vec_out <= "1000111101011011011111111011110101011001111110111111000100100010";
                    when "01011" => level_vec_out <= "1000111101011011011111111011110101011001111110111111000100100010";
                    when "01100" => level_vec_out <= "1000111101011011011111111011110101011001111110111111000100100010";
                    when "01101" => level_vec_out <= "1001111101011011011111111011110101011001111110111111000100100010";
                    when "01110" => level_vec_out <= "1001111101011011111111111011110101011001111110111111000100100010";
                    when "01111" => level_vec_out <= "1001111101011011111111111011111101011101111110111111000100100010";
                    when "10000" => level_vec_out <= "1001111101011011111111111011111101011101111110111111000110100010";
                    when "10001" => level_vec_out <= "1001111101011011111111111011111101011101111111111111000110110010";
                    when "10010" => level_vec_out <= "1001111101011011111111111011111101011101111111111111000110110010";
                    when "10011" => level_vec_out <= "1001111111011011111111111011111101011101111111111111000110110010";
                    when "10100" => level_vec_out <= "1011111111011011111111111011111111011101111111111111000110110010";
                    when "10101" => level_vec_out <= "1011111111111011111111111111111111011101111111111111001110110010";
                    when "10110" => level_vec_out <= "1011111111111011111111111111111111011101111111111111001110110010";
                    when "10111" => level_vec_out <= "1111111111111011111111111111111111011101111111111111001111110010";
                    when "11000" => level_vec_out <= "1111111111111011111111111111111111111101111111111111001111110010";
                    when "11001" => level_vec_out <= "1111111111111011111111111111111111111101111111111111001111110011";
                    when "11010" => level_vec_out <= "1111111111111011111111111111111111111111111111111111001111110011";
                    when "11011" => level_vec_out <= "1111111111111011111111111111111111111111111111111111011111110011";
                    when "11100" => level_vec_out <= "1111111111111011111111111111111111111111111111111111011111110011";
                    when "11101" => level_vec_out <= "1111111111111111111111111111111111111111111111111111011111110011";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111111111111111011111110111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "001" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0110001110010010100111110111010100110001011110111101110110011001";
                    when "00001" => level_vec_out <= "1110001110010111100111110111010100110001011110111101110110011001";
                    when "00010" => level_vec_out <= "1110001110010111100111110111010100110001011110111101110110011001";
                    when "00011" => level_vec_out <= "1110001110010111100111110111010100110001111110111101110110011001";
                    when "00100" => level_vec_out <= "1110001111010111100111110111010110110001111110111101110110011001";
                    when "00101" => level_vec_out <= "1110001111010111100111110111010110110001111110111101110110011001";
                    when "00110" => level_vec_out <= "1110001111010111100111110111010110111101111110111101110110011001";
                    when "00111" => level_vec_out <= "1110001111010111110111110111010110111101111110111101110110011001";
                    when "01000" => level_vec_out <= "1110001111010111110111110111010110111101111110111101110110011001";
                    when "01001" => level_vec_out <= "1110001111010111110111110111010110111101111110111101110110011001";
                    when "01010" => level_vec_out <= "1111001111010111110111110111010110111101111110111101110110011001";
                    when "01011" => level_vec_out <= "1111001111010111110111110111010110111101111110111101110110011001";
                    when "01100" => level_vec_out <= "1111001111010111110111110111010110111101111110111101110110111001";
                    when "01101" => level_vec_out <= "1111001111010111110111110111110110111101111110111101110110111001";
                    when "01110" => level_vec_out <= "1111001111010111110111110111111110111101111110111111110110111101";
                    when "01111" => level_vec_out <= "1111001111010111110111110111111110111101111110111111110110111101";
                    when "10000" => level_vec_out <= "1111001111010111110111110111111110111101111110111111110110111101";
                    when "10001" => level_vec_out <= "1111001111010111110111110111111110111101111110111111110110111101";
                    when "10010" => level_vec_out <= "1111001111010111110111110111111110111101111110111111110110111101";
                    when "10011" => level_vec_out <= "1111001111010111110111110111111110111101111110111111110110111101";
                    when "10100" => level_vec_out <= "1111001111010111110111111111111110111101111110111111110110111101";
                    when "10101" => level_vec_out <= "1111011111010111110111111111111110111111111111111111110110111101";
                    when "10110" => level_vec_out <= "1111011111010111111111111111111110111111111111111111111110111101";
                    when "10111" => level_vec_out <= "1111011111010111111111111111111110111111111111111111111110111101";
                    when "11000" => level_vec_out <= "1111011111010111111111111111111110111111111111111111111111111101";
                    when "11001" => level_vec_out <= "1111011111010111111111111111111110111111111111111111111111111101";
                    when "11010" => level_vec_out <= "1111111111010111111111111111111110111111111111111111111111111101";
                    when "11011" => level_vec_out <= "1111111111010111111111111111111110111111111111111111111111111111";
                    when "11100" => level_vec_out <= "1111111111010111111111111111111111111111111111111111111111111111";
                    when "11101" => level_vec_out <= "1111111111010111111111111111111111111111111111111111111111111111";
                    when "11110" => level_vec_out <= "1111111111011111111111111111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "010" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1011001101100100100001001011100111000111011000000011001011110101";
                    when "00001" => level_vec_out <= "1011001101100100100001001011100111000111011000000011001011110101";
                    when "00010" => level_vec_out <= "1011001101100100100001001011100111000111011101000011001011110101";
                    when "00011" => level_vec_out <= "1011001101100100100001001011100111000111011101000011001011110101";
                    when "00100" => level_vec_out <= "1011001101100100100001001011100111000111011101000011001011110101";
                    when "00101" => level_vec_out <= "1011001101100100100001001011100111000111011101000011001011110101";
                    when "00110" => level_vec_out <= "1011001101100100100001001011100111000111011101010011001011110101";
                    when "00111" => level_vec_out <= "1011001101100100100001001011100111000111011101010011001011111101";
                    when "01000" => level_vec_out <= "1011001101100100100011001011101111000111011101010011001111111101";
                    when "01001" => level_vec_out <= "1011001101100100100011001011101111001111011101010011001111111101";
                    when "01010" => level_vec_out <= "1011001101100100100011001011101111001111011101010011001111111101";
                    when "01011" => level_vec_out <= "1011001101100100100011001011101111001111111101010011001111111101";
                    when "01100" => level_vec_out <= "1011001101100100100011001011101111001111111101011011001111111101";
                    when "01101" => level_vec_out <= "1011001101101100110011001011101111001111111101011011001111111101";
                    when "01110" => level_vec_out <= "1011001101101100110011001011101111001111111101011011001111111101";
                    when "01111" => level_vec_out <= "1011001101101100110011011011101111001111111101111011001111111101";
                    when "10000" => level_vec_out <= "1111001101101100110111011011101111001111111101111011001111111101";
                    when "10001" => level_vec_out <= "1111001101101110110111011011101111001111111101111011001111111101";
                    when "10010" => level_vec_out <= "1111001101101110110111011011101111011111111111111011101111111101";
                    when "10011" => level_vec_out <= "1111001101101110110111011011101111011111111111111011101111111101";
                    when "10100" => level_vec_out <= "1111001101101110110111011011111111011111111111111011101111111101";
                    when "10101" => level_vec_out <= "1111001101101110110111011011111111011111111111111011101111111101";
                    when "10110" => level_vec_out <= "1111001101101110110111011011111111011111111111111011101111111101";
                    when "10111" => level_vec_out <= "1111001101101111110111011011111111011111111111111011101111111101";
                    when "11000" => level_vec_out <= "1111001101101111110111111011111111011111111111111011101111111101";
                    when "11001" => level_vec_out <= "1111001101111111110111111011111111111111111111111011101111111101";
                    when "11010" => level_vec_out <= "1111001101111111110111111011111111111111111111111011101111111101";
                    when "11011" => level_vec_out <= "1111001111111111110111111011111111111111111111111011101111111111";
                    when "11100" => level_vec_out <= "1111001111111111110111111111111111111111111111111011111111111111";
                    when "11101" => level_vec_out <= "1111001111111111110111111111111111111111111111111011111111111111";
                    when "11110" => level_vec_out <= "1111001111111111111111111111111111111111111111111011111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111011111111111111";
                when others => null;
                end case;
            when "011" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0101000010011011010111110101010001111000111000101010101101100111";
                    when "00001" => level_vec_out <= "0101000010011011010111110101010001111000111000101010101101100111";
                    when "00010" => level_vec_out <= "0101000110011011010111110101010001111000111000101010101101101111";
                    when "00011" => level_vec_out <= "1111000110011011010111111101010001111000111000101010101101101111";
                    when "00100" => level_vec_out <= "1111000110011011010111111101010001111000111000101110101101101111";
                    when "00101" => level_vec_out <= "1111000110011011010111111101110101111000111000101110101101101111";
                    when "00110" => level_vec_out <= "1111000110011011010111111101110101111000111000101110101111101111";
                    when "00111" => level_vec_out <= "1111000110011011010111111101110101111000111000101110101111101111";
                    when "01000" => level_vec_out <= "1111001110011011010111111101111101111000111000101110101111111111";
                    when "01001" => level_vec_out <= "1111001110011011011111111101111101111000111000101110101111111111";
                    when "01010" => level_vec_out <= "1111011110011011111111111101111101111000111000101110101111111111";
                    when "01011" => level_vec_out <= "1111011110011011111111111101111101111000111100101110101111111111";
                    when "01100" => level_vec_out <= "1111011110011011111111111101111101111000111100101110101111111111";
                    when "01101" => level_vec_out <= "1111011110011011111111111111111101111000111100101110101111111111";
                    when "01110" => level_vec_out <= "1111011111011011111111111111111101111000111100101110101111111111";
                    when "01111" => level_vec_out <= "1111011111011011111111111111111111111000111100101110101111111111";
                    when "10000" => level_vec_out <= "1111011111011011111111111111111111111000111101101110101111111111";
                    when "10001" => level_vec_out <= "1111011111011011111111111111111111111000111101101110101111111111";
                    when "10010" => level_vec_out <= "1111011111011011111111111111111111111000111111111110101111111111";
                    when "10011" => level_vec_out <= "1111011111011011111111111111111111111000111111111110101111111111";
                    when "10100" => level_vec_out <= "1111011111011011111111111111111111111000111111111110101111111111";
                    when "10101" => level_vec_out <= "1111011111011011111111111111111111111000111111111110101111111111";
                    when "10110" => level_vec_out <= "1111011111011011111111111111111111111000111111111110101111111111";
                    when "10111" => level_vec_out <= "1111011111111011111111111111111111111000111111111110101111111111";
                    when "11000" => level_vec_out <= "1111111111111011111111111111111111111000111111111110101111111111";
                    when "11001" => level_vec_out <= "1111111111111011111111111111111111111000111111111110101111111111";
                    when "11010" => level_vec_out <= "1111111111111111111111111111111111111100111111111110101111111111";
                    when "11011" => level_vec_out <= "1111111111111111111111111111111111111100111111111110101111111111";
                    when "11100" => level_vec_out <= "1111111111111111111111111111111111111100111111111111111111111111";
                    when "11101" => level_vec_out <= "1111111111111111111111111111111111111101111111111111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111101111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111101111111111111111111111111";
                when others => null;
                end case;
            when "100" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0000000101111001000100001011010001110111010001000100100110110010";
                    when "00001" => level_vec_out <= "0000000101111001000100001011010001110111010001000100100110110010";
                    when "00010" => level_vec_out <= "0000000101111001000100001011010001110111010001000100100110110010";
                    when "00011" => level_vec_out <= "0000000101111001000100001011010001110111010001000100100110110010";
                    when "00100" => level_vec_out <= "0000000101111001000100001011010001110111010001000100111110110010";
                    when "00101" => level_vec_out <= "0000000101111001000100001111010001110111010001000100111110110010";
                    when "00110" => level_vec_out <= "0000000101111001000100001111010001110111010001000100111110110110";
                    when "00111" => level_vec_out <= "0000000101111001001100101111010001110111010001000100111110110110";
                    when "01000" => level_vec_out <= "0000000101111001001100101111010001110111010001000100111110110110";
                    when "01001" => level_vec_out <= "0000000101111001001100101111010001110111010001000100111111110111";
                    when "01010" => level_vec_out <= "0000000101111001001100101111010001110111010001100100111111110111";
                    when "01011" => level_vec_out <= "0000000101111011001100101111010001110111010001100100111111111111";
                    when "01100" => level_vec_out <= "0000000101111011001100101111011001110111010001100100111111111111";
                    when "01101" => level_vec_out <= "0000000101111011001100101111011001110111010001100100111111111111";
                    when "01110" => level_vec_out <= "0000000101111011001100101111011011110111010001100100111111111111";
                    when "01111" => level_vec_out <= "0000000101111011001100101111011011110111010001100101111111111111";
                    when "10000" => level_vec_out <= "0001001101111111001100101111011011110111011001100101111111111111";
                    when "10001" => level_vec_out <= "0001001101111111011100101111011011110111111001100101111111111111";
                    when "10010" => level_vec_out <= "0011001101111111011100101111011011110111111001100101111111111111";
                    when "10011" => level_vec_out <= "0011001111111111011100101111011011110111111011100101111111111111";
                    when "10100" => level_vec_out <= "0111001111111111011100101111111011110111111011100101111111111111";
                    when "10101" => level_vec_out <= "0111001111111111011100101111111011110111111011110101111111111111";
                    when "10110" => level_vec_out <= "1111001111111111011101101111111011110111111011110101111111111111";
                    when "10111" => level_vec_out <= "1111011111111111011101101111111111110111111011110101111111111111";
                    when "11000" => level_vec_out <= "1111011111111111011101101111111111111111111011110101111111111111";
                    when "11001" => level_vec_out <= "1111011111111111011101101111111111111111111011110101111111111111";
                    when "11010" => level_vec_out <= "1111011111111111011101101111111111111111111011110101111111111111";
                    when "11011" => level_vec_out <= "1111011111111111011101111111111111111111111011110101111111111111";
                    when "11100" => level_vec_out <= "1111111111111111011101111111111111111111111011110101111111111111";
                    when "11101" => level_vec_out <= "1111111111111111011101111111111111111111111111110101111111111111";
                    when "11110" => level_vec_out <= "1111111111111111011101111111111111111111111111110111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111101111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "101" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0100101110101000011000010010000101010011010001000110000110001000";
                    when "00001" => level_vec_out <= "0100101110101000011000010010000101010011010001000110000110001000";
                    when "00010" => level_vec_out <= "0100101110101000011000010010100101011011010001000110000110001000";
                    when "00011" => level_vec_out <= "0100111110111000011000010010100101011011010001000110000110001000";
                    when "00100" => level_vec_out <= "0100111110111000011000010010100101011011010001000110000110001000";
                    when "00101" => level_vec_out <= "0100111110111000011010010010100101011011010001000110000110101000";
                    when "00110" => level_vec_out <= "0100111110111000011010010010100101011011010001000110000110101000";
                    when "00111" => level_vec_out <= "0100111110111000011010110010100101011111010001000110000110101000";
                    when "01000" => level_vec_out <= "0100111110111000011010110010100101011111010001000110000110101000";
                    when "01001" => level_vec_out <= "0100111110111001011010110010100101011111010001100110010110101000";
                    when "01010" => level_vec_out <= "0110111110111001011010110011100101011111011001100110010110101000";
                    when "01011" => level_vec_out <= "0110111110111001011110110011100101011111011001100110010110101000";
                    when "01100" => level_vec_out <= "0110111110111001011110110011100101011111011101100111010110101000";
                    when "01101" => level_vec_out <= "0110111110111001011110110011100101011111011101100111010111111000";
                    when "01110" => level_vec_out <= "0110111110111001011110110011100101011111011101100111010111111000";
                    when "01111" => level_vec_out <= "0110111110111001011110110011100101011111011101100111010111111000";
                    when "10000" => level_vec_out <= "0110111110111001011110110011100101011111011101100111010111111000";
                    when "10001" => level_vec_out <= "0110111110111001011110110011101101011111011101110111010111111001";
                    when "10010" => level_vec_out <= "0111111110111001011110110011101101011111011101110111010111111001";
                    when "10011" => level_vec_out <= "0111111110111011011110110011111101011111011101110111110111111001";
                    when "10100" => level_vec_out <= "0111111110111011011110110011111101011111011101110111110111111001";
                    when "10101" => level_vec_out <= "0111111110111011011110111011111101011111011101110111110111111001";
                    when "10110" => level_vec_out <= "0111111110111111011110111011111101111111111101110111110111111001";
                    when "10111" => level_vec_out <= "0111111110111111011110111011111101111111111111110111110111111001";
                    when "11000" => level_vec_out <= "0111111110111111011110111011111101111111111111110111110111111001";
                    when "11001" => level_vec_out <= "0111111110111111011110111011111101111111111111110111110111111011";
                    when "11010" => level_vec_out <= "0111111110111111011110111011111101111111111111110111110111111011";
                    when "11011" => level_vec_out <= "0111111110111111011111111011111101111111111111110111110111111011";
                    when "11100" => level_vec_out <= "0111111110111111011111111011111101111111111111110111110111111111";
                    when "11101" => level_vec_out <= "0111111110111111111111111011111101111111111111110111110111111111";
                    when "11110" => level_vec_out <= "1111111110111111111111111011111111111111111111111111110111111111";
                    when "11111" => level_vec_out <= "1111111110111111111111111011111111111111111111111111110111111111";
                when others => null;
                end case;
            when "110" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1110011111000100001001011111001001111101110011000110101001001101";
                    when "00001" => level_vec_out <= "1110011111000100001011011111001001111111110011000110101001001101";
                    when "00010" => level_vec_out <= "1110011111000100001011011111001001111111110011000110101001001101";
                    when "00011" => level_vec_out <= "1110011111000100001011011111001011111111110011000110101001001101";
                    when "00100" => level_vec_out <= "1110011111000100001011011111001011111111110011000110101001001101";
                    when "00101" => level_vec_out <= "1111011111100100001011011111001011111111110011000110101001001101";
                    when "00110" => level_vec_out <= "1111011111100100001011011111001011111111110011100110101001001101";
                    when "00111" => level_vec_out <= "1111011111100100001011011111001011111111110011100110101001001101";
                    when "01000" => level_vec_out <= "1111011111100100011111011111001011111111110011100110101001001101";
                    when "01001" => level_vec_out <= "1111011111100100111111011111001011111111110011100110101001001101";
                    when "01010" => level_vec_out <= "1111011111100100111111011111001011111111110011100110101001001101";
                    when "01011" => level_vec_out <= "1111011111100100111111011111011011111111110011100111101001011101";
                    when "01100" => level_vec_out <= "1111011111101100111111011111011011111111110011100111101101011101";
                    when "01101" => level_vec_out <= "1111011111101110111111011111011011111111110011100111101101011101";
                    when "01110" => level_vec_out <= "1111011111101110111111011111011011111111111011100111101101011101";
                    when "01111" => level_vec_out <= "1111011111101110111111011111011011111111111011100111101111011101";
                    when "10000" => level_vec_out <= "1111011111101110111111011111011011111111111011100111101111011101";
                    when "10001" => level_vec_out <= "1111011111101110111111011111011011111111111011100111101111011101";
                    when "10010" => level_vec_out <= "1111011111101110111111011111111011111111111011100111101111011101";
                    when "10011" => level_vec_out <= "1111011111101110111111011111111011111111111011110111101111011101";
                    when "10100" => level_vec_out <= "1111111111101110111111011111111111111111111011110111101111011101";
                    when "10101" => level_vec_out <= "1111111111101110111111011111111111111111111011110111101111011101";
                    when "10110" => level_vec_out <= "1111111111101110111111011111111111111111111011110111101111011101";
                    when "10111" => level_vec_out <= "1111111111101110111111011111111111111111111011110111101111011101";
                    when "11000" => level_vec_out <= "1111111111101110111111011111111111111111111011111111111111011101";
                    when "11001" => level_vec_out <= "1111111111111111111111011111111111111111111011111111111111011101";
                    when "11010" => level_vec_out <= "1111111111111111111111011111111111111111111011111111111111111101";
                    when "11011" => level_vec_out <= "1111111111111111111111011111111111111111111011111111111111111101";
                    when "11100" => level_vec_out <= "1111111111111111111111011111111111111111111011111111111111111101";
                    when "11101" => level_vec_out <= "1111111111111111111111111111111111111111111011111111111111111101";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111111011111111111111111101";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111011111111111111111101";
                when others => null;
                end case;
            when "111" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0101111110111110010111011011111110010010011011101000001111111001";
                    when "00001" => level_vec_out <= "0101111110111110010111011011111110110010011011101000001111111001";
                    when "00010" => level_vec_out <= "0101111110111110010111011011111110110010011011101000001111111001";
                    when "00011" => level_vec_out <= "0101111110111110010111011011111110110010011011101000001111111001";
                    when "00100" => level_vec_out <= "0101111110111110010111011011111110110010011111101000001111111001";
                    when "00101" => level_vec_out <= "0101111110111110010111011011111110110010011111101000001111111001";
                    when "00110" => level_vec_out <= "0101111110111110010111011011111110110010011111101000001111111001";
                    when "00111" => level_vec_out <= "0101111110111110010111011011111110110010011111101000001111111001";
                    when "01000" => level_vec_out <= "0101111110111110010111011011111110110010011111101000001111111001";
                    when "01001" => level_vec_out <= "0101111110111110010111011011111110110010011111101000001111111001";
                    when "01010" => level_vec_out <= "0101111110111110010111011011111110110010011111101001001111111001";
                    when "01011" => level_vec_out <= "0101111110111110010111011011111110110010011111101001001111111001";
                    when "01100" => level_vec_out <= "0101111110111110010111011011111110110010111111101001001111111001";
                    when "01101" => level_vec_out <= "0101111110111110010111011011111110110010111111101001001111111001";
                    when "01110" => level_vec_out <= "1101111110111110010111011011111110110010111111101001001111111001";
                    when "01111" => level_vec_out <= "1101111110111110010111011011111110110010111111101101001111111001";
                    when "10000" => level_vec_out <= "1101111110111110010111011011111110110010111111101101001111111001";
                    when "10001" => level_vec_out <= "1101111110111110010111011011111110110010111111101101001111111001";
                    when "10010" => level_vec_out <= "1101111110111110010111011011111110110010111111101101001111111001";
                    when "10011" => level_vec_out <= "1101111110111110011111011011111110110010111111101101001111111001";
                    when "10100" => level_vec_out <= "1101111110111110011111011011111110110010111111101101001111111001";
                    when "10101" => level_vec_out <= "1101111110111110011111011011111110110010111111101101001111111001";
                    when "10110" => level_vec_out <= "1101111110111110011111111011111110110010111111101101001111111001";
                    when "10111" => level_vec_out <= "1101111110111110011111111011111110110010111111101101001111111101";
                    when "11000" => level_vec_out <= "1101111110111110011111111011111110110010111111111101001111111101";
                    when "11001" => level_vec_out <= "1101111110111110011111111011111110110110111111111101011111111101";
                    when "11010" => level_vec_out <= "1101111110111110111111111111111110111110111111111101011111111101";
                    when "11011" => level_vec_out <= "1111111110111110111111111111111110111110111111111101011111111111";
                    when "11100" => level_vec_out <= "1111111110111110111111111111111110111111111111111101011111111111";
                    when "11101" => level_vec_out <= "1111111111111110111111111111111111111111111111111101111111111111";
                    when "11110" => level_vec_out <= "1111111111111110111111111111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when others => null;
        end case;
    end process;
end Behavioral;