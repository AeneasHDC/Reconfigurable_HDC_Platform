----
 -- @file level_hvec_gen_hdl.hpp
 -- @brief This script generates HDL code for generating high-dimensional LEVEL vectors.
 -- It is a novel method; for more information, please refer to our paper.
 --
 -- @author Saeid Jamili and Marco Angioli
 -- @note Author names are listed in alphabetical order.
 -- @email <saeid.jamili@uniroma1.it>
 -- @email <marco.angioli@uniroma1.it>
 --
 -- @contributors
 --
 -- @date Created: 24th July 2023
 -- @date Last Updated: 23th August 2023
 --
 -- @version 1.0.0
 --
 -- @institute Sapienza University of Rome
 -- @cite https://doi.org/10.xxxx/yyyyy
 --
 -- @section DEPENDENCIES
 -- - Dependency1: Description or version details.
 -- - Dependency2: Description or version details.
 --
 -- @section LICENSE
 -- This file is part of the Aeneas HyperCompute Platform.
 --
 -- Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 --
 -- @section CHANGELOG
 -- @version 1.0.0-dev - 23th August 2023
 -- - Initial release
 --
 -- @todo
 -- - Complete level vector generator function
 -- - Add training
 --
 -- @see
 -- -
 -- -
 -- -
 --
 --

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity level_vec_gen is
    Port ( level_vec_out : out  STD_LOGIC_VECTOR (63 downto 0);
           frame_index : in  STD_LOGIC_VECTOR (2 downto 0);
           frame_id : in  STD_LOGIC_VECTOR (4 downto 0));
end level_vec_gen;

architecture Behavioral of level_vec_gen is
begin
    process (frame_index, frame_id)
    begin
        -- Update this function to match your requirements
        case frame_index is
            when "000" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0001000101000110010001011010001110011011100010011011000100101100";
                    when "00001" => level_vec_out <= "0001000101000110010001011010001110011011100010011011000100101100";
                    when "00010" => level_vec_out <= "0001000101000110010001011010001110011011100010011011000101101100";
                    when "00011" => level_vec_out <= "0001000101000110010001011010001110011011100010011011000101101100";
                    when "00100" => level_vec_out <= "0001000101000110010001011010001110011011100010011011000101101100";
                    when "00101" => level_vec_out <= "0001000101000110010001011010001110011011100010011011000101101100";
                    when "00110" => level_vec_out <= "0001000101000110010001011110001110011011100110011011000101101100";
                    when "00111" => level_vec_out <= "0001000101000110010001011110001110011011100110011111000101101100";
                    when "01000" => level_vec_out <= "0001010101000110010001011110001110011011100110011111000101101100";
                    when "01001" => level_vec_out <= "0001010101000110010001111110001110011011100110011111000101101100";
                    when "01010" => level_vec_out <= "0011010101000110010001111110001110011011100110011111000101101100";
                    when "01011" => level_vec_out <= "0011110101000110010001111110001110011011100110011111010101101100";
                    when "01100" => level_vec_out <= "1011110101000110010011111110101110011011100110011111010101101100";
                    when "01101" => level_vec_out <= "1011110101000110010011111110101110011011101110011111010101101100";
                    when "01110" => level_vec_out <= "1011110101000110010011111110101110011011101110011111010101101100";
                    when "01111" => level_vec_out <= "1011110101000110010011111110101110011011101110011111011101101100";
                    when "10000" => level_vec_out <= "1011110101000110010011111110101110011011101110011111011101101100";
                    when "10001" => level_vec_out <= "1011110101000110010011111110101110011011101110011111011101101100";
                    when "10010" => level_vec_out <= "1011111101010110010011111110101110011011111110011111011101101100";
                    when "10011" => level_vec_out <= "1011111101010110010011111110111110011011111111011111111101101100";
                    when "10100" => level_vec_out <= "1011111101010110010011111110111111011011111111011111111101101110";
                    when "10101" => level_vec_out <= "1011111101010110010011111110111111011011111111011111111101101110";
                    when "10110" => level_vec_out <= "1011111101010110010111111111111111011011111111011111111111101110";
                    when "10111" => level_vec_out <= "1011111101010110010111111111111111011011111111011111111111101110";
                    when "11000" => level_vec_out <= "1011111101110110010111111111111111011011111111011111111111101110";
                    when "11001" => level_vec_out <= "1011111111110110111111111111111111011111111111011111111111101110";
                    when "11010" => level_vec_out <= "1011111111111110111111111111111111011111111111011111111111101110";
                    when "11011" => level_vec_out <= "1011111111111110111111111111111111011111111111011111111111101111";
                    when "11100" => level_vec_out <= "1011111111111110111111111111111111111111111111011111111111101111";
                    when "11101" => level_vec_out <= "1011111111111110111111111111111111111111111111011111111111101111";
                    when "11110" => level_vec_out <= "1111111111111110111111111111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111110111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "001" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0111000000100110000111011100111011001011101110101001011111000110";
                    when "00001" => level_vec_out <= "0111000000100110000111011101111011001011101110101001011111000110";
                    when "00010" => level_vec_out <= "0111000000100110000111011101111011001011111110101001011111000110";
                    when "00011" => level_vec_out <= "0111000000100110000111011101111011001011111111101001011111000110";
                    when "00100" => level_vec_out <= "0111000000100110000111011101111011001011111111101011011111000111";
                    when "00101" => level_vec_out <= "0111000000100110000111011101111011001011111111101011011111000111";
                    when "00110" => level_vec_out <= "0111000001100110000111011101111011001011111111101011011111000111";
                    when "00111" => level_vec_out <= "0111000001100110000111011101111011001011111111101111011111000111";
                    when "01000" => level_vec_out <= "0111000001100111000111011101111011001011111111101111011111000111";
                    when "01001" => level_vec_out <= "1111000001101111000111011101111011001011111111101111011111000111";
                    when "01010" => level_vec_out <= "1111000011101111000111011101111011001011111111101111011111000111";
                    when "01011" => level_vec_out <= "1111000011101111000111011101111011001011111111101111011111000111";
                    when "01100" => level_vec_out <= "1111000011101111000111011101111011001011111111101111011111000111";
                    when "01101" => level_vec_out <= "1111000011101111000111011101111011001011111111101111011111000111";
                    when "01110" => level_vec_out <= "1111000011101111000111011101111111001011111111101111011111000111";
                    when "01111" => level_vec_out <= "1111001011101111000111011101111111001011111111101111011111000111";
                    when "10000" => level_vec_out <= "1111001111101111100111011111111111001011111111101111011111000111";
                    when "10001" => level_vec_out <= "1111001111101111100111011111111111001111111111101111011111100111";
                    when "10010" => level_vec_out <= "1111001111101111100111011111111111001111111111101111011111100111";
                    when "10011" => level_vec_out <= "1111011111101111110111011111111111001111111111101111011111100111";
                    when "10100" => level_vec_out <= "1111011111101111110111011111111111011111111111101111011111100111";
                    when "10101" => level_vec_out <= "1111011111101111111111011111111111011111111111111111011111100111";
                    when "10110" => level_vec_out <= "1111011111111111111111011111111111011111111111111111011111100111";
                    when "10111" => level_vec_out <= "1111011111111111111111011111111111011111111111111111111111100111";
                    when "11000" => level_vec_out <= "1111011111111111111111011111111111011111111111111111111111100111";
                    when "11001" => level_vec_out <= "1111011111111111111111011111111111011111111111111111111111110111";
                    when "11010" => level_vec_out <= "1111011111111111111111011111111111011111111111111111111111110111";
                    when "11011" => level_vec_out <= "1111011111111111111111111111111111011111111111111111111111110111";
                    when "11100" => level_vec_out <= "1111011111111111111111111111111111011111111111111111111111111111";
                    when "11101" => level_vec_out <= "1111111111111111111111111111111111011111111111111111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111011111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111011111111111111111111111111111";
                when others => null;
                end case;
            when "010" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0110011011111111100011110001100111100001101110111011001110111010";
                    when "00001" => level_vec_out <= "0110011011111111100011110001100111100001101110111011001110111010";
                    when "00010" => level_vec_out <= "0110011011111111100011110101100111100001101110111011001110111010";
                    when "00011" => level_vec_out <= "0110011011111111100011110101100111100001111110111011001110111010";
                    when "00100" => level_vec_out <= "0110011011111111100011110101100111100001111110111011001110111010";
                    when "00101" => level_vec_out <= "0110011011111111100011110111100111100001111110111011001110111010";
                    when "00110" => level_vec_out <= "0110011011111111100011110111100111100001111110111011001110111110";
                    when "00111" => level_vec_out <= "0110111011111111100011110111100111100001111110111011001110111110";
                    when "01000" => level_vec_out <= "0110111011111111100011111111100111100001111110111011001110111110";
                    when "01001" => level_vec_out <= "0110111011111111100011111111110111100001111110111011001110111110";
                    when "01010" => level_vec_out <= "0110111011111111100011111111110111100101111110111011001111111110";
                    when "01011" => level_vec_out <= "0110111011111111100011111111110111100101111110111011011111111110";
                    when "01100" => level_vec_out <= "0110111011111111100011111111110111100101111110111011011111111110";
                    when "01101" => level_vec_out <= "0110111011111111100011111111110111100101111110111011011111111110";
                    when "01110" => level_vec_out <= "0110111011111111110011111111110111100101111110111011011111111110";
                    when "01111" => level_vec_out <= "0110111111111111111011111111110111100101111110111011011111111110";
                    when "10000" => level_vec_out <= "0110111111111111111011111111110111100101111110111011011111111110";
                    when "10001" => level_vec_out <= "0110111111111111111011111111110111100101111110111011011111111110";
                    when "10010" => level_vec_out <= "0110111111111111111011111111110111100101111110111011011111111110";
                    when "10011" => level_vec_out <= "0110111111111111111011111111110111100101111110111011011111111110";
                    when "10100" => level_vec_out <= "0110111111111111111011111111110111101101111110111011011111111110";
                    when "10101" => level_vec_out <= "0110111111111111111011111111110111101101111110111011011111111110";
                    when "10110" => level_vec_out <= "0110111111111111111011111111110111101101111110111011011111111111";
                    when "10111" => level_vec_out <= "1110111111111111111011111111110111101101111110111011011111111111";
                    when "11000" => level_vec_out <= "1110111111111111111011111111110111111101111110111011011111111111";
                    when "11001" => level_vec_out <= "1110111111111111111111111111110111111101111110111011011111111111";
                    when "11010" => level_vec_out <= "1110111111111111111111111111111111111101111110111011011111111111";
                    when "11011" => level_vec_out <= "1110111111111111111111111111111111111101111111111111011111111111";
                    when "11100" => level_vec_out <= "1110111111111111111111111111111111111101111111111111011111111111";
                    when "11101" => level_vec_out <= "1110111111111111111111111111111111111101111111111111011111111111";
                    when "11110" => level_vec_out <= "1110111111111111111111111111111111111101111111111111011111111111";
                    when "11111" => level_vec_out <= "1110111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "011" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1100101111100000101011110110010001101000110000000011000111110001";
                    when "00001" => level_vec_out <= "1110101111100000101011110110010001101000110000000011000111110001";
                    when "00010" => level_vec_out <= "1110101111100000101011110110010001101000110100000011000111110001";
                    when "00011" => level_vec_out <= "1111101111100000101011110110010001101000110100000111000111110011";
                    when "00100" => level_vec_out <= "1111101111100000101011110110110001101000110100010111000111110011";
                    when "00101" => level_vec_out <= "1111101111100100101011110110110001101000110101010111000111110011";
                    when "00110" => level_vec_out <= "1111101111100100101011110110110001111000110101010111000111110011";
                    when "00111" => level_vec_out <= "1111101111100100101011110110110001111000110101110111000111110011";
                    when "01000" => level_vec_out <= "1111101111100100101111111110110001111000110101110111000111110011";
                    when "01001" => level_vec_out <= "1111101111100100101111111110110001111000110101111111000111110011";
                    when "01010" => level_vec_out <= "1111101111100100101111111111110001111000110101111111001111110011";
                    when "01011" => level_vec_out <= "1111101111110100101111111111110001111000110101111111001111110011";
                    when "01100" => level_vec_out <= "1111101111110100101111111111110001111000110111111111001111110011";
                    when "01101" => level_vec_out <= "1111101111110100101111111111110001111001110111111111001111110011";
                    when "01110" => level_vec_out <= "1111101111110110101111111111110001111001110111111111001111110011";
                    when "01111" => level_vec_out <= "1111101111110110101111111111110001111001110111111111001111110011";
                    when "10000" => level_vec_out <= "1111101111110110101111111111110001111001110111111111001111110011";
                    when "10001" => level_vec_out <= "1111101111110110101111111111110001111001110111111111001111110011";
                    when "10010" => level_vec_out <= "1111101111110110101111111111110101111001110111111111001111110011";
                    when "10011" => level_vec_out <= "1111101111110110101111111111110101111001110111111111001111110011";
                    when "10100" => level_vec_out <= "1111101111110110101111111111110101111001110111111111001111110011";
                    when "10101" => level_vec_out <= "1111101111110110101111111111110101111001110111111111001111110011";
                    when "10110" => level_vec_out <= "1111101111110110111111111111111101111001110111111111001111110011";
                    when "10111" => level_vec_out <= "1111101111111110111111111111111101111001110111111111001111110011";
                    when "11000" => level_vec_out <= "1111101111111110111111111111111101111001110111111111011111110111";
                    when "11001" => level_vec_out <= "1111101111111110111111111111111101111001110111111111011111110111";
                    when "11010" => level_vec_out <= "1111101111111110111111111111111101111011110111111111011111111111";
                    when "11011" => level_vec_out <= "1111101111111110111111111111111101111011110111111111011111111111";
                    when "11100" => level_vec_out <= "1111111111111110111111111111111101111011110111111111011111111111";
                    when "11101" => level_vec_out <= "1111111111111111111111111111111101111011110111111111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111101111011110111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111101111111111111111111111111111111";
                when others => null;
                end case;
            when "100" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0001110111100001011100101100010000011010001000001000001000111100";
                    when "00001" => level_vec_out <= "0001110111100001011100101100010000011111001000001000001100111100";
                    when "00010" => level_vec_out <= "0001110111100001011100101100110000011111001000001000001100111100";
                    when "00011" => level_vec_out <= "0001110111100001111100101100110000011111001000001000001100111100";
                    when "00100" => level_vec_out <= "0001110111100001111100101100110000011111001100001001001100111100";
                    when "00101" => level_vec_out <= "0001110111100001111100101100110000011111001110011001001100111100";
                    when "00110" => level_vec_out <= "0001110111100001111100101100111000011111001110011001011100111100";
                    when "00111" => level_vec_out <= "0001110111100001111100101100111000011111001110011001111100111100";
                    when "01000" => level_vec_out <= "0001110111100001111100101100111000011111001110011001111100111100";
                    when "01001" => level_vec_out <= "0001110111100001111100101100111000011111001110011001111100111100";
                    when "01010" => level_vec_out <= "0001110111100001111100101100111000011111001110011001111100111100";
                    when "01011" => level_vec_out <= "0001110111100001111100101100111000011111001110011011111100111110";
                    when "01100" => level_vec_out <= "0001111111100001111100101100111000111111001110011011111100111111";
                    when "01101" => level_vec_out <= "0001111111100001111110101100111000111111001110011011111100111111";
                    when "01110" => level_vec_out <= "0001111111100001111110101100111000111111001110011011111100111111";
                    when "01111" => level_vec_out <= "0001111111100001111110101100111000111111001110111011111100111111";
                    when "10000" => level_vec_out <= "0001111111100001111110101100111001111111011110111011111100111111";
                    when "10001" => level_vec_out <= "0001111111100001111111111100111001111111011110111011111100111111";
                    when "10010" => level_vec_out <= "0001111111100001111111111100111001111111011110111011111100111111";
                    when "10011" => level_vec_out <= "0001111111100001111111111100111001111111011110111011111100111111";
                    when "10100" => level_vec_out <= "0001111111100101111111111100111001111111011110111011111100111111";
                    when "10101" => level_vec_out <= "0011111111110101111111111101111001111111011110111111111100111111";
                    when "10110" => level_vec_out <= "0011111111110101111111111101111001111111011110111111111100111111";
                    when "10111" => level_vec_out <= "0011111111110111111111111101111001111111011110111111111100111111";
                    when "11000" => level_vec_out <= "0011111111110111111111111101111101111111011110111111111100111111";
                    when "11001" => level_vec_out <= "0011111111110111111111111101111101111111011110111111111100111111";
                    when "11010" => level_vec_out <= "0011111111110111111111111101111101111111011110111111111100111111";
                    when "11011" => level_vec_out <= "0011111111110111111111111101111101111111011110111111111110111111";
                    when "11100" => level_vec_out <= "0011111111110111111111111101111101111111011111111111111110111111";
                    when "11101" => level_vec_out <= "0111111111110111111111111101111101111111011111111111111110111111";
                    when "11110" => level_vec_out <= "1111111111110111111111111101111101111111011111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111101111111011111111111111111111111";
                when others => null;
                end case;
            when "101" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0001100101001100101000000000111001100010000110110011101110001011";
                    when "00001" => level_vec_out <= "0001100101001110101000000000111001100010000110110011111110001011";
                    when "00010" => level_vec_out <= "1001101101001110101000000000111001100010000110110011111110001011";
                    when "00011" => level_vec_out <= "1001101101001110101000000000111001100010000110110011111110001011";
                    when "00100" => level_vec_out <= "1001101101001110101000000010111001100010000110110011111110001011";
                    when "00101" => level_vec_out <= "1001101101001110101000010010111001100010000110110011111110101011";
                    when "00110" => level_vec_out <= "1001101101001110101000010010111001100010000110111011111110101011";
                    when "00111" => level_vec_out <= "1001101101001110111000010010111001100010000110111011111110101011";
                    when "01000" => level_vec_out <= "1001101101001110111000010010111001100010000110111011111110101011";
                    when "01001" => level_vec_out <= "1001101101001110111000010010111001100010000110111011111110101011";
                    when "01010" => level_vec_out <= "1001101101011110111000010010111001100010000110111011111110101011";
                    when "01011" => level_vec_out <= "1001101101011110111000010010111001100010010110111011111110101011";
                    when "01100" => level_vec_out <= "1001101101011110111000010010111001100010010110111011111110101011";
                    when "01101" => level_vec_out <= "1001101101011110111001010010111001100010010110111011111110101111";
                    when "01110" => level_vec_out <= "1001101101011110111001011010111001100110010110111011111110101111";
                    when "01111" => level_vec_out <= "1001101101011111111001011010111001100110010110111011111110101111";
                    when "10000" => level_vec_out <= "1001101101011111111001011010111001100110010111111011111110101111";
                    when "10001" => level_vec_out <= "1001101101011111111001011010111001100111010111111111111110101111";
                    when "10010" => level_vec_out <= "1011101101011111111001011010111101100111010111111111111110101111";
                    when "10011" => level_vec_out <= "1011101101011111111011011010111101100111010111111111111110101111";
                    when "10100" => level_vec_out <= "1011101101011111111011011010111101100111110111111111111110101111";
                    when "10101" => level_vec_out <= "1011101101011111111011011010111101100111110111111111111110101111";
                    when "10110" => level_vec_out <= "1011101101011111111011011010111101100111110111111111111110101111";
                    when "10111" => level_vec_out <= "1011101101011111111111111010111101101111110111111111111111101111";
                    when "11000" => level_vec_out <= "1011101101011111111111111110111101101111111111111111111111101111";
                    when "11001" => level_vec_out <= "1011101101011111111111111110111101101111111111111111111111101111";
                    when "11010" => level_vec_out <= "1011101101011111111111111110111101111111111111111111111111101111";
                    when "11011" => level_vec_out <= "1011101101011111111111111110111101111111111111111111111111101111";
                    when "11100" => level_vec_out <= "1011111101011111111111111110111101111111111111111111111111111111";
                    when "11101" => level_vec_out <= "1011111111011111111111111110111101111111111111111111111111111111";
                    when "11110" => level_vec_out <= "1111111111011111111111111110111101111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111101111111111111111111111111111111";
                when others => null;
                end case;
            when "110" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0010010101100101010110110110111011000111010011000111101010011111";
                    when "00001" => level_vec_out <= "0011010101100101010110110110111011000111010011000111101010011111";
                    when "00010" => level_vec_out <= "0011010101100101010110110111111011000111010011000111101010011111";
                    when "00011" => level_vec_out <= "0011010101100101010110110111111011000111011011000111101010011111";
                    when "00100" => level_vec_out <= "0011010101100111010110110111111011000111011011000111101010011111";
                    when "00101" => level_vec_out <= "0011010101100111010110110111111011000111011011000111101010011111";
                    when "00110" => level_vec_out <= "0011010101100111010110110111111011000111011011000111101010011111";
                    when "00111" => level_vec_out <= "0011010101100111010110110111111011000111011011000111101010011111";
                    when "01000" => level_vec_out <= "0011010101100111010110110111111011000111011011000111101010111111";
                    when "01001" => level_vec_out <= "0011010101100111011110110111111011000111011011000111101010111111";
                    when "01010" => level_vec_out <= "0011010101100111011110110111111011000111011011000111101110111111";
                    when "01011" => level_vec_out <= "0011010101100111011110110111111011000111011011010111101110111111";
                    when "01100" => level_vec_out <= "0011010101100111011110110111111011000111011011010111101110111111";
                    when "01101" => level_vec_out <= "0111110101100111011110110111111011000111011011010111111110111111";
                    when "01110" => level_vec_out <= "0111110101100111011110110111111011100111011111010111111110111111";
                    when "01111" => level_vec_out <= "1111110101100111011110110111111011100111011111010111111110111111";
                    when "10000" => level_vec_out <= "1111110101100111011110110111111011110111011111010111111110111111";
                    when "10001" => level_vec_out <= "1111110101100111011110110111111011110111111111010111111110111111";
                    when "10010" => level_vec_out <= "1111111101100111011110111111111011110111111111010111111110111111";
                    when "10011" => level_vec_out <= "1111111101100111011110111111111111110111111111010111111110111111";
                    when "10100" => level_vec_out <= "1111111101100111011110111111111111111111111111010111111111111111";
                    when "10101" => level_vec_out <= "1111111101100111011110111111111111111111111111010111111111111111";
                    when "10110" => level_vec_out <= "1111111101100111011110111111111111111111111111010111111111111111";
                    when "10111" => level_vec_out <= "1111111101100111011110111111111111111111111111010111111111111111";
                    when "11000" => level_vec_out <= "1111111101100111011110111111111111111111111111010111111111111111";
                    when "11001" => level_vec_out <= "1111111101100111011110111111111111111111111111010111111111111111";
                    when "11010" => level_vec_out <= "1111111101100111011110111111111111111111111111111111111111111111";
                    when "11011" => level_vec_out <= "1111111111110111111110111111111111111111111111111111111111111111";
                    when "11100" => level_vec_out <= "1111111111110111111110111111111111111111111111111111111111111111";
                    when "11101" => level_vec_out <= "1111111111111111111110111111111111111111111111111111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "111" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1011001011011010111010010011111011000110111001111110110011000100";
                    when "00001" => level_vec_out <= "1011001011011010111010010011111011000110111001111110110011000100";
                    when "00010" => level_vec_out <= "1011001011011010111010010011111011000110111001111110110011000100";
                    when "00011" => level_vec_out <= "1011001011111010111010010011111011000110111001111110110011000100";
                    when "00100" => level_vec_out <= "1011001011111010111010010011111011000110111001111110110011000100";
                    when "00101" => level_vec_out <= "1011001011111010111010110011111011000110111001111110110011000100";
                    when "00110" => level_vec_out <= "1011001011111010111010110011111011000110111001111110110011000100";
                    when "00111" => level_vec_out <= "1011001111111010111011110011111011000110111001111110110011000100";
                    when "01000" => level_vec_out <= "1011001111111011111011110011111011000110111011111110110011000100";
                    when "01001" => level_vec_out <= "1011001111111011111011110011111111000110111011111111110011000100";
                    when "01010" => level_vec_out <= "1011001111111011111011110011111111000110111011111111110011000100";
                    when "01011" => level_vec_out <= "1011001111111011111011110011111111000110111011111111110011000100";
                    when "01100" => level_vec_out <= "1011001111111011111011110011111111000110111111111111110011000100";
                    when "01101" => level_vec_out <= "1011001111111011111011110011111111000110111111111111110011000100";
                    when "01110" => level_vec_out <= "1011001111111011111011110011111111000110111111111111110011000101";
                    when "01111" => level_vec_out <= "1011001111111011111011110011111111000110111111111111110011100101";
                    when "10000" => level_vec_out <= "1011001111111011111011110011111111010110111111111111110011100101";
                    when "10001" => level_vec_out <= "1011001111111011111011110011111111010110111111111111111011100101";
                    when "10010" => level_vec_out <= "1011001111111011111011110011111111010110111111111111111011100101";
                    when "10011" => level_vec_out <= "1011001111111111111011110011111111010110111111111111111011100101";
                    when "10100" => level_vec_out <= "1011001111111111111011110011111111010110111111111111111011100101";
                    when "10101" => level_vec_out <= "1011001111111111111011111011111111011110111111111111111011100101";
                    when "10110" => level_vec_out <= "1011001111111111111011111011111111011111111111111111111011100101";
                    when "10111" => level_vec_out <= "1011001111111111111011111011111111011111111111111111111011100101";
                    when "11000" => level_vec_out <= "1011001111111111111011111011111111011111111111111111111111100101";
                    when "11001" => level_vec_out <= "1011001111111111111011111111111111111111111111111111111111100101";
                    when "11010" => level_vec_out <= "1011001111111111111111111111111111111111111111111111111111100101";
                    when "11011" => level_vec_out <= "1011001111111111111111111111111111111111111111111111111111100101";
                    when "11100" => level_vec_out <= "1111001111111111111111111111111111111111111111111111111111110101";
                    when "11101" => level_vec_out <= "1111011111111111111111111111111111111111111111111111111111111101";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111101";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111101";
                when others => null;
                end case;
            when others => null;
        end case;
    end process;
end Behavioral;