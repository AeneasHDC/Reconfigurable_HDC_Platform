/**
 * @file level_hvec_gen_hdl.hpp
 * @brief This script generates HDL code for generating high-dimensional LEVEL vectors.
 * It is a novel method; for more information, please refer to our paper.
 *
 * @author Saeid Jamili and Marco Angioli
 * @note Author names are listed in alphabetical order.
 * @email <saeid.jamili@uniroma1.it>
 * @email <marco.angioli@uniroma1.it>
 *
 * @contributors
 *
 * @date Created: 24th July 2023
 * @date Last Updated: 23th August 2023
 *
 * @version 1.0.0
 *
 * @institute Sapienza University of Rome
 * @cite https://doi.org/10.xxxx/yyyyy
 *
 * @section DEPENDENCIES
 * - Dependency1: Description or version details.
 * - Dependency2: Description or version details.
 *
 * @section LICENSE
 * This file is part of the Aeneas HyperCompute Platform.
 *
 * Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 *
 * @section CHANGELOG
 * @version 1.0.0-dev - 23th August 2023
 * - Initial release
 *
 * @todo
 * - Complete level vector generator function
 * - Add training
 *
 * @see
 * -
 * -
 * -
 *
 */

module level_hvec_gen #(parameter int DI_PARALLEL_W_BITS = 64) (
  input logic [2:0] frame_index,
  input logic [4:0] frame_id,
  output logic [DI_PARALLEL_W_BITS-1:0] level_vec_out
);
  always_comb begin
    case (frame_index)
      0:
        case (frame_id)
          0:
            level_vec_out = 64'b1110101001000111011010001101101011111000010001010010011000100100;
          1:
            level_vec_out = 64'b1110101001000111011010001101101011111000010001010010011000100100;
          2:
            level_vec_out = 64'b1110101001000111011010001101101011111000010001010010011000100100;
          3:
            level_vec_out = 64'b1110101001000111011010001101101011111010010001010010011000100100;
          4:
            level_vec_out = 64'b1110101001010111011010101101101011111010010001010010011000101100;
          5:
            level_vec_out = 64'b1110101001010111011010101101101011111010010001010010011000101110;
          6:
            level_vec_out = 64'b1110101001011111011010101101101011111010010001011010011000101110;
          7:
            level_vec_out = 64'b1110101001011111011010101101101011111010010001011010011000101110;
          8:
            level_vec_out = 64'b1110101001011111011010101101101011111010010001011010011000101110;
          9:
            level_vec_out = 64'b1110101001011111011010101101101011111110010001011010111000101110;
          10:
            level_vec_out = 64'b1110101101011111011010111101101011111111010001011110111000101110;
          11:
            level_vec_out = 64'b1110101101011111011010111101101011111111010001011110111000101110;
          12:
            level_vec_out = 64'b1110101101011111011010111111101011111111010001011110111000101110;
          13:
            level_vec_out = 64'b1111101101011111011010111111101011111111010001011110111000101110;
          14:
            level_vec_out = 64'b1111101101011111111010111111101011111111110001011111111000101110;
          15:
            level_vec_out = 64'b1111101101011111111010111111101011111111110001011111111000101110;
          16:
            level_vec_out = 64'b1111101101011111111010111111111011111111111001011111111000101110;
          17:
            level_vec_out = 64'b1111101101011111111010111111111011111111111001011111111001101110;
          18:
            level_vec_out = 64'b1111101101011111111010111111111011111111111001011111111001101110;
          19:
            level_vec_out = 64'b1111101101011111111010111111111011111111111001011111111001101110;
          20:
            level_vec_out = 64'b1111101101011111111010111111111111111111111001011111111001101110;
          21:
            level_vec_out = 64'b1111101101011111111010111111111111111111111001111111111001101110;
          22:
            level_vec_out = 64'b1111101101011111111010111111111111111111111001111111111001101110;
          23:
            level_vec_out = 64'b1111101101011111111110111111111111111111111001111111111001101110;
          24:
            level_vec_out = 64'b1111101101011111111110111111111111111111111001111111111001101110;
          25:
            level_vec_out = 64'b1111101111011111111110111111111111111111111001111111111001101110;
          26:
            level_vec_out = 64'b1111101111011111111110111111111111111111111101111111111001101110;
          27:
            level_vec_out = 64'b1111101111011111111110111111111111111111111101111111111101101110;
          28:
            level_vec_out = 64'b1111101111011111111111111111111111111111111101111111111101101110;
          29:
            level_vec_out = 64'b1111101111011111111111111111111111111111111101111111111101111110;
          30:
            level_vec_out = 64'b1111111111011111111111111111111111111111111101111111111101111111;
          31:
            level_vec_out = 64'b1111111111011111111111111111111111111111111111111111111101111111;
        endcase
      1:
        case (frame_id)
          0:
            level_vec_out = 64'b0010100001011000000101101000010011110110100011000100111110100010;
          1:
            level_vec_out = 64'b0010100001011000000101101000010011110110100011000100111110100010;
          2:
            level_vec_out = 64'b0010111001111000000101101000010011110110100011000100111110100010;
          3:
            level_vec_out = 64'b0010111101111000000101101000010011110110100011000100111110100010;
          4:
            level_vec_out = 64'b0010111101111000000101101000010011110110100011000100111110100010;
          5:
            level_vec_out = 64'b0011111101111000000101101000010011110110110011000100111110100110;
          6:
            level_vec_out = 64'b0011111101111000000101101000010011110110110111010110111110100110;
          7:
            level_vec_out = 64'b0011111101111000000101101000110111110110110111010110111110100110;
          8:
            level_vec_out = 64'b0011111101111000000101101000110111110110110111010110111110100110;
          9:
            level_vec_out = 64'b0011111101111000000101101100110111110110110111010110111110100110;
          10:
            level_vec_out = 64'b0011111101111000000101101100110111110110110111010110111110100110;
          11:
            level_vec_out = 64'b1011111101111000001101101100110111110110110111010110111110100110;
          12:
            level_vec_out = 64'b1011111101111000001101101100110111110110110111110110111110110110;
          13:
            level_vec_out = 64'b1011111101111000001101101100110111110110110111110110111110110110;
          14:
            level_vec_out = 64'b1011111101111010001101101100110111110110110111110110111110110110;
          15:
            level_vec_out = 64'b1011111101111010011101101100110111110110110111110110111110110111;
          16:
            level_vec_out = 64'b1011111101111010011101101110110111110110110111110110111111110111;
          17:
            level_vec_out = 64'b1011111111111010011101101110110111110110110111110110111111110111;
          18:
            level_vec_out = 64'b1011111111111010011101101110110111110110111111110111111111110111;
          19:
            level_vec_out = 64'b1011111111111010011111101110110111110110111111110111111111110111;
          20:
            level_vec_out = 64'b1011111111111010011111101110110111111110111111110111111111110111;
          21:
            level_vec_out = 64'b1011111111111010011111101110111111111110111111110111111111110111;
          22:
            level_vec_out = 64'b1011111111111010111111101110111111111110111111110111111111110111;
          23:
            level_vec_out = 64'b1011111111111010111111101110111111111110111111110111111111110111;
          24:
            level_vec_out = 64'b1011111111111011111111101110111111111110111111110111111111110111;
          25:
            level_vec_out = 64'b1011111111111011111111101110111111111110111111110111111111110111;
          26:
            level_vec_out = 64'b1011111111111011111111101110111111111110111111110111111111110111;
          27:
            level_vec_out = 64'b1011111111111011111111101111111111111110111111111111111111110111;
          28:
            level_vec_out = 64'b1011111111111111111111101111111111111110111111111111111111110111;
          29:
            level_vec_out = 64'b1011111111111111111111101111111111111110111111111111111111111111;
          30:
            level_vec_out = 64'b1011111111111111111111101111111111111111111111111111111111111111;
          31:
            level_vec_out = 64'b1111111111111111111111101111111111111111111111111111111111111111;
        endcase
      2:
        case (frame_id)
          0:
            level_vec_out = 64'b1101100111011100001000001001010000010101100010010111001000010111;
          1:
            level_vec_out = 64'b1101100111011100001000001001010000010101100010010111001000010111;
          2:
            level_vec_out = 64'b1101100111011100001000001001010000010101100010010111001000010111;
          3:
            level_vec_out = 64'b1101100111011100001000001001010001011101100010010111001000010111;
          4:
            level_vec_out = 64'b1101100111011100001000001001010001011101100010010111001000110111;
          5:
            level_vec_out = 64'b1101100111011100001000001001010001011101100010010111011000110111;
          6:
            level_vec_out = 64'b1101100111011100001010001001010001011101100010010111011000110111;
          7:
            level_vec_out = 64'b1101100111011101001010001001010001011101100010010111011000110111;
          8:
            level_vec_out = 64'b1101100111011101001010001101010001011111100010010111011000110111;
          9:
            level_vec_out = 64'b1101100111011101101010001101010001011111100010010111011000110111;
          10:
            level_vec_out = 64'b1101100111011101101010001101010001011111100010010111011000110111;
          11:
            level_vec_out = 64'b1101100111011101101010001101010001011111100010010111011000110111;
          12:
            level_vec_out = 64'b1101100111011101101010001101010001011111100010010111011001110111;
          13:
            level_vec_out = 64'b1101100111011101101010001101010001011111100010010111011001110111;
          14:
            level_vec_out = 64'b1101100111011101101010001101011001011111100010110111011001110111;
          15:
            level_vec_out = 64'b1101100111011101101010001101011001011111100010110111011001110111;
          16:
            level_vec_out = 64'b1101100111011101101010001101011001111111100010111111011001110111;
          17:
            level_vec_out = 64'b1101100111011101101010001101011101111111100010111111011001110111;
          18:
            level_vec_out = 64'b1101100111011111101010001101011101111111100010111111011001110111;
          19:
            level_vec_out = 64'b1101100111011111101010001101011101111111100010111111011001110111;
          20:
            level_vec_out = 64'b1101100111011111101010001101011101111111100010111111011101110111;
          21:
            level_vec_out = 64'b1101101111011111101010001101011101111111100010111111011101110111;
          22:
            level_vec_out = 64'b1101101111011111111010001101011111111111100011111111111101110111;
          23:
            level_vec_out = 64'b1101101111111111111010001101011111111111100011111111111101110111;
          24:
            level_vec_out = 64'b1101101111111111111011001101011111111111110011111111111111110111;
          25:
            level_vec_out = 64'b1101101111111111111011001101011111111111110011111111111111111111;
          26:
            level_vec_out = 64'b1101101111111111111011001101011111111111111011111111111111111111;
          27:
            level_vec_out = 64'b1111101111111111111011001101011111111111111011111111111111111111;
          28:
            level_vec_out = 64'b1111101111111111111011001111011111111111111011111111111111111111;
          29:
            level_vec_out = 64'b1111101111111111111011001111111111111111111111111111111111111111;
          30:
            level_vec_out = 64'b1111101111111111111111101111111111111111111111111111111111111111;
          31:
            level_vec_out = 64'b1111101111111111111111111111111111111111111111111111111111111111;
        endcase
      3:
        case (frame_id)
          0:
            level_vec_out = 64'b1011000101111000101000111010111011110101001000011110011111011111;
          1:
            level_vec_out = 64'b1011000101111000101000111110111011110101001000011110011111011111;
          2:
            level_vec_out = 64'b1011000101111000101000111110111011110101001000011110011111011111;
          3:
            level_vec_out = 64'b1011000101111000101000111110111011110101001000011110011111011111;
          4:
            level_vec_out = 64'b1011001101111000111000111110111011110101001000011110011111011111;
          5:
            level_vec_out = 64'b1011001101111000111000111110111011110101001000011110011111011111;
          6:
            level_vec_out = 64'b1011001101111000111000111110111011110101001000011110011111011111;
          7:
            level_vec_out = 64'b1011001101111000111000111110111011110101001000011110011111011111;
          8:
            level_vec_out = 64'b1011101101111000111000111110111011110101001000011111011111011111;
          9:
            level_vec_out = 64'b1011101101111100111000111110111011110101001000011111011111011111;
          10:
            level_vec_out = 64'b1011101101111100111000111110111011110101001000011111011111011111;
          11:
            level_vec_out = 64'b1011101101111100111000111110111011110101001010011111011111011111;
          12:
            level_vec_out = 64'b1011111101111100111000111110111011110101001010011111011111011111;
          13:
            level_vec_out = 64'b1111111101111101111000111110111011110101001010011111011111011111;
          14:
            level_vec_out = 64'b1111111101111101111000111110111011110101001110011111011111011111;
          15:
            level_vec_out = 64'b1111111101111101111000111110111011110101001110111111011111011111;
          16:
            level_vec_out = 64'b1111111101111101111010111110111011110101001110111111011111011111;
          17:
            level_vec_out = 64'b1111111101111101111010111110111011110101101110111111011111111111;
          18:
            level_vec_out = 64'b1111111101111101111010111110111011110101101110111111111111111111;
          19:
            level_vec_out = 64'b1111111101111101111010111110111011110111101110111111111111111111;
          20:
            level_vec_out = 64'b1111111101111101111010111110111011110111101110111111111111111111;
          21:
            level_vec_out = 64'b1111111101111101111010111110111011110111101111111111111111111111;
          22:
            level_vec_out = 64'b1111111101111111111010111110111011110111101111111111111111111111;
          23:
            level_vec_out = 64'b1111111101111111111010111110111011110111101111111111111111111111;
          24:
            level_vec_out = 64'b1111111101111111111010111110111011111111111111111111111111111111;
          25:
            level_vec_out = 64'b1111111101111111111010111110111011111111111111111111111111111111;
          26:
            level_vec_out = 64'b1111111101111111111110111110111111111111111111111111111111111111;
          27:
            level_vec_out = 64'b1111111101111111111110111110111111111111111111111111111111111111;
          28:
            level_vec_out = 64'b1111111111111111111110111110111111111111111111111111111111111111;
          29:
            level_vec_out = 64'b1111111111111111111110111110111111111111111111111111111111111111;
          30:
            level_vec_out = 64'b1111111111111111111110111110111111111111111111111111111111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111110111111111111111111111111111111111111;
        endcase
      4:
        case (frame_id)
          0:
            level_vec_out = 64'b1100011101010000111000011110001111010010000101001010110110111000;
          1:
            level_vec_out = 64'b1100011101010000111000011110001111010010000101001010110110111101;
          2:
            level_vec_out = 64'b1100011101010000111000011110011111010010000101001010110110111101;
          3:
            level_vec_out = 64'b1100011101010000111000011110011111010010000101001010110110111101;
          4:
            level_vec_out = 64'b1100011101010000111000011111011111010010000101001010110110111101;
          5:
            level_vec_out = 64'b1100011101010000111000011111011111010010000101001010110110111101;
          6:
            level_vec_out = 64'b1100011101010000111000011111011111010010000101001010110110111101;
          7:
            level_vec_out = 64'b1100011101010000111000011111011111010010000101101010110111111101;
          8:
            level_vec_out = 64'b1100011101010000111000011111011111010010000101101010110111111101;
          9:
            level_vec_out = 64'b1100011101010000111000011111011111010010000101101010110111111101;
          10:
            level_vec_out = 64'b1100011101010000111000111111011111010010000101101010110111111101;
          11:
            level_vec_out = 64'b1100011101011000111000111111011111010010000101101110111111111101;
          12:
            level_vec_out = 64'b1110011101011000111000111111011111010010000101101110111111111101;
          13:
            level_vec_out = 64'b1110011101011000111000111111011111110010000101101110111111111101;
          14:
            level_vec_out = 64'b1110011101011000111000111111011111110010000101101110111111111101;
          15:
            level_vec_out = 64'b1110011101011000111000111111011111110010000101101110111111111101;
          16:
            level_vec_out = 64'b1110011101011000111000111111011111110010000101101110111111111101;
          17:
            level_vec_out = 64'b1110011101011000111000111111011111110010000101101110111111111101;
          18:
            level_vec_out = 64'b1110011101011000111000111111011111110010000101111110111111111101;
          19:
            level_vec_out = 64'b1110011101111000111000111111111111110010000101111110111111111111;
          20:
            level_vec_out = 64'b1110011101111000111010111111111111110010010101111110111111111111;
          21:
            level_vec_out = 64'b1110011101111000111010111111111111110010010101111110111111111111;
          22:
            level_vec_out = 64'b1110111101111010111010111111111111110010010101111110111111111111;
          23:
            level_vec_out = 64'b1110111101111010111010111111111111110011010111111110111111111111;
          24:
            level_vec_out = 64'b1110111101111010111010111111111111110011010111111110111111111111;
          25:
            level_vec_out = 64'b1110111111111011111010111111111111110011010111111110111111111111;
          26:
            level_vec_out = 64'b1110111111111011111110111111111111110011010111111110111111111111;
          27:
            level_vec_out = 64'b1110111111111011111110111111111111110111010111111110111111111111;
          28:
            level_vec_out = 64'b1111111111111011111110111111111111110111010111111110111111111111;
          29:
            level_vec_out = 64'b1111111111111011111110111111111111110111010111111111111111111111;
          30:
            level_vec_out = 64'b1111111111111111111110111111111111110111011111111111111111111111;
          31:
            level_vec_out = 64'b1111111111111111111110111111111111110111111111111111111111111111;
        endcase
      5:
        case (frame_id)
          0:
            level_vec_out = 64'b1101110001101000001100011110000101110101101011010001011101001001;
          1:
            level_vec_out = 64'b1101110001101000001100011110000101110101101011010001011101001011;
          2:
            level_vec_out = 64'b1101110001101000001100011110000101110101101011010001011101001011;
          3:
            level_vec_out = 64'b1101110001101000001100011110000101110101101011010001011101001011;
          4:
            level_vec_out = 64'b1101110001101000001100011110000101110101101011010001011101001011;
          5:
            level_vec_out = 64'b1101110001101000011100011110000101110101101011010001011101011011;
          6:
            level_vec_out = 64'b1101110001101000011100011110000101110101101011010001011101011011;
          7:
            level_vec_out = 64'b1101110001101000011100011110010101110101101011010001011101011011;
          8:
            level_vec_out = 64'b1101110001101100011100011110010101110101101011010001011101011011;
          9:
            level_vec_out = 64'b1101110001101100011100011110010101110111101011010001011101011011;
          10:
            level_vec_out = 64'b1111110001101100011101011110110101110111101011010001011101011011;
          11:
            level_vec_out = 64'b1111110001101100011101011110110101110111101011010001011101011011;
          12:
            level_vec_out = 64'b1111110001101100011101011110110101110111101011010001011101011111;
          13:
            level_vec_out = 64'b1111110001101100011101011110111101110111101011010001011101011111;
          14:
            level_vec_out = 64'b1111110001101100011101011110111101110111101011010001011101011111;
          15:
            level_vec_out = 64'b1111110001101100011101011110111101110111101011011001011101011111;
          16:
            level_vec_out = 64'b1111110001101100011101011110111101110111101011011001011101011111;
          17:
            level_vec_out = 64'b1111111001101101011101011110111101110111101011011101011101011111;
          18:
            level_vec_out = 64'b1111111001111101011101011110111101110111101011011111011101011111;
          19:
            level_vec_out = 64'b1111111001111101011101011110111101110111101011011111111101011111;
          20:
            level_vec_out = 64'b1111111001111101011101011111111101111111101011011111111101011111;
          21:
            level_vec_out = 64'b1111111001111101011101011111111101111111101011011111111111011111;
          22:
            level_vec_out = 64'b1111111001111101011101011111111101111111101011011111111111011111;
          23:
            level_vec_out = 64'b1111111001111101011101011111111101111111111011011111111111011111;
          24:
            level_vec_out = 64'b1111111001111101011101011111111101111111111011011111111111011111;
          25:
            level_vec_out = 64'b1111111001111111011101011111111101111111111111011111111111011111;
          26:
            level_vec_out = 64'b1111111101111111011101011111111111111111111111011111111111011111;
          27:
            level_vec_out = 64'b1111111101111111111101011111111111111111111111011111111111011111;
          28:
            level_vec_out = 64'b1111111101111111111101011111111111111111111111011111111111111111;
          29:
            level_vec_out = 64'b1111111111111111111101011111111111111111111111011111111111111111;
          30:
            level_vec_out = 64'b1111111111111111111111011111111111111111111111011111111111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111011111111111111111;
        endcase
      6:
        case (frame_id)
          0:
            level_vec_out = 64'b1111111101100011010101000001110110010001010011100100000110101001;
          1:
            level_vec_out = 64'b1111111101100011110101000001110110010011010011100100010110101001;
          2:
            level_vec_out = 64'b1111111101100011110101000011110110010011010011100100010110101001;
          3:
            level_vec_out = 64'b1111111101100011110101010011110110010011111011100100010110101001;
          4:
            level_vec_out = 64'b1111111101100011110101010011110110010011111011100100010110101001;
          5:
            level_vec_out = 64'b1111111101100011110101010011110110010011111011100100010110101001;
          6:
            level_vec_out = 64'b1111111101100011110101010111110110010011111011100100010110101001;
          7:
            level_vec_out = 64'b1111111101100011110101010111110110010011111011100100010110101101;
          8:
            level_vec_out = 64'b1111111101100011111101010111111110010011111011100100010110101101;
          9:
            level_vec_out = 64'b1111111101100011111101010111111110011011111011110100010110101101;
          10:
            level_vec_out = 64'b1111111101100011111101010111111110011011111011110100010110101101;
          11:
            level_vec_out = 64'b1111111101100011111101010111111110111011111011110100010110111101;
          12:
            level_vec_out = 64'b1111111101100011111101010111111110111011111011110100010110111101;
          13:
            level_vec_out = 64'b1111111101100111111101110111111110111011111011110100010110111101;
          14:
            level_vec_out = 64'b1111111101101111111101110111111110111011111011110100010110111101;
          15:
            level_vec_out = 64'b1111111101101111111101110111111110111011111011110100010110111101;
          16:
            level_vec_out = 64'b1111111101101111111101111111111110111011111011110100010110111101;
          17:
            level_vec_out = 64'b1111111101101111111101111111111110111011111011110100010110111101;
          18:
            level_vec_out = 64'b1111111101101111111101111111111110111011111011110110010110111101;
          19:
            level_vec_out = 64'b1111111101101111111101111111111110111011111011110111010110111101;
          20:
            level_vec_out = 64'b1111111101101111111101111111111110111011111011110111010110111101;
          21:
            level_vec_out = 64'b1111111101101111111111111111111110111011111011110111110111111101;
          22:
            level_vec_out = 64'b1111111101101111111111111111111110111011111011110111110111111101;
          23:
            level_vec_out = 64'b1111111101101111111111111111111110111111111011110111110111111101;
          24:
            level_vec_out = 64'b1111111101101111111111111111111110111111111011110111110111111101;
          25:
            level_vec_out = 64'b1111111111101111111111111111111110111111111011110111110111111101;
          26:
            level_vec_out = 64'b1111111111101111111111111111111111111111111011110111110111111101;
          27:
            level_vec_out = 64'b1111111111101111111111111111111111111111111011110111110111111111;
          28:
            level_vec_out = 64'b1111111111111111111111111111111111111111111011110111110111111111;
          29:
            level_vec_out = 64'b1111111111111111111111111111111111111111111011111111111111111111;
          30:
            level_vec_out = 64'b1111111111111111111111111111111111111111111011111111111111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        endcase
      7:
        case (frame_id)
          0:
            level_vec_out = 64'b0100001111011001111011111100100000111101101101111010101101010011;
          1:
            level_vec_out = 64'b0100001111011001111011111100101000111101101101111010101101010011;
          2:
            level_vec_out = 64'b0100011111011001111011111100101000111111111101111010101101010011;
          3:
            level_vec_out = 64'b0100011111011001111011111100101000111111111101111010101111010011;
          4:
            level_vec_out = 64'b0100011111111001111011111100101000111111111101111010101111010011;
          5:
            level_vec_out = 64'b0100011111111001111011111100101000111111111101111110101111010011;
          6:
            level_vec_out = 64'b0100011111111001111011111100111000111111111101111110101111010011;
          7:
            level_vec_out = 64'b0100011111111001111011111100111001111111111101111110101111010011;
          8:
            level_vec_out = 64'b0100111111111001111011111100111001111111111101111110101111010011;
          9:
            level_vec_out = 64'b0100111111111001111011111100111001111111111101111110101111010011;
          10:
            level_vec_out = 64'b0100111111111001111011111100111001111111111101111110101111010011;
          11:
            level_vec_out = 64'b0100111111111001111011111100111001111111111101111110101111010011;
          12:
            level_vec_out = 64'b0100111111111001111111111100111001111111111101111110101111010011;
          13:
            level_vec_out = 64'b0100111111111011111111111100111001111111111101111110101111010011;
          14:
            level_vec_out = 64'b0100111111111011111111111100111001111111111101111110101111010011;
          15:
            level_vec_out = 64'b1100111111111011111111111110111001111111111101111110111111011011;
          16:
            level_vec_out = 64'b1100111111111011111111111110111001111111111101111110111111011011;
          17:
            level_vec_out = 64'b1100111111111011111111111110111001111111111101111110111111011011;
          18:
            level_vec_out = 64'b1100111111111011111111111110111001111111111101111110111111011011;
          19:
            level_vec_out = 64'b1110111111111011111111111110111001111111111101111110111111011011;
          20:
            level_vec_out = 64'b1110111111111111111111111110111001111111111101111110111111011011;
          21:
            level_vec_out = 64'b1110111111111111111111111110111001111111111101111110111111011011;
          22:
            level_vec_out = 64'b1110111111111111111111111110111001111111111101111110111111011011;
          23:
            level_vec_out = 64'b1110111111111111111111111110111101111111111101111110111111011111;
          24:
            level_vec_out = 64'b1110111111111111111111111111111111111111111101111110111111011111;
          25:
            level_vec_out = 64'b1111111111111111111111111111111111111111111101111110111111011111;
          26:
            level_vec_out = 64'b1111111111111111111111111111111111111111111101111110111111011111;
          27:
            level_vec_out = 64'b1111111111111111111111111111111111111111111101111110111111111111;
          28:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111110111111111111;
          29:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111110111111111111;
          30:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111110111111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        endcase
    endcase
  end
endmodule