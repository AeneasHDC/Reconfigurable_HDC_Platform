/**
 * @file level_hvec_gen_hdl.hpp
 * @brief This script generates HDL code for generating high-dimensional LEVEL vectors.
 * It is a novel method; for more information, please refer to our paper.
 *
 * @author Saeid Jamili and Marco Angioli
 * @note Author names are listed in alphabetical order.
 * @email <saeid.jamili@uniroma1.it>
 * @email <marco.angioli@uniroma1.it>
 *
 * @contributors
 *
 * @date Created: 24th July 2023
 * @date Last Updated: 23th August 2023
 *
 * @version 1.0.0
 *
 * @institute Sapienza University of Rome
 * @cite https://doi.org/10.xxxx/yyyyy
 *
 * @section DEPENDENCIES
 * - Dependency1: Description or version details.
 * - Dependency2: Description or version details.
 *
 * @section LICENSE
 * This file is part of the Aeneas HyperCompute Platform.
 *
 * Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 *
 * @section CHANGELOG
 * @version 1.0.0-dev - 23th August 2023
 * - Initial release
 *
 * @todo
 * - Complete level vector generator function
 * - Add training
 *
 * @see
 * -
 * -
 * -
 *
 */

module level_hvec_gen #(parameter int DI_PARALLEL_W_BITS = 64) (
  input logic [2:0] frame_index,
  input logic [4:0] frame_id,
  output logic [DI_PARALLEL_W_BITS-1:0] level_vec_out
);
  always_comb begin
    case (frame_index)
      0:
        case (frame_id)
          0:
            level_vec_out = 64'b0110101000011000111110101101110110100100010101110101000000111111;
          1:
            level_vec_out = 64'b0110101000011000111110101101110110100100010101110101000000111111;
          2:
            level_vec_out = 64'b0110111000011000111110101101110110100100010101110101100001111111;
          3:
            level_vec_out = 64'b0110111101011000111110101101110110100100010101110101100001111111;
          4:
            level_vec_out = 64'b0110111101011000111110101101110110100100010101110101100001111111;
          5:
            level_vec_out = 64'b1110111101011000111110101101110110100100010101110101100001111111;
          6:
            level_vec_out = 64'b1110111101011000111110101101110110100100010101110101100001111111;
          7:
            level_vec_out = 64'b1110111111011000111111101101110110101100010101110101100001111111;
          8:
            level_vec_out = 64'b1110111111011000111111101101110110101100010101110101100001111111;
          9:
            level_vec_out = 64'b1110111111011000111111101101110110101100010101110101101001111111;
          10:
            level_vec_out = 64'b1110111111011000111111101101110110101100010101110101101001111111;
          11:
            level_vec_out = 64'b1110111111011010111111101101110110101100011101110101101001111111;
          12:
            level_vec_out = 64'b1110111111011010111111101101110110101100011101111101101001111111;
          13:
            level_vec_out = 64'b1110111111011010111111101101110110101100011101111101111001111111;
          14:
            level_vec_out = 64'b1110111111011010111111101101110110101100011101111101111001111111;
          15:
            level_vec_out = 64'b1110111111011110111111101101110110101100011111111101111001111111;
          16:
            level_vec_out = 64'b1110111111011110111111111101110110101100011111111101111001111111;
          17:
            level_vec_out = 64'b1111111111011110111111111101110110101100011111111101111001111111;
          18:
            level_vec_out = 64'b1111111111011110111111111101110110101100011111111111111001111111;
          19:
            level_vec_out = 64'b1111111111011110111111111101110110101100011111111111111001111111;
          20:
            level_vec_out = 64'b1111111111011110111111111101110110101110011111111111111001111111;
          21:
            level_vec_out = 64'b1111111111011110111111111101110110101110011111111111111001111111;
          22:
            level_vec_out = 64'b1111111111011110111111111101110111101110011111111111111001111111;
          23:
            level_vec_out = 64'b1111111111011110111111111101110111101111011111111111111001111111;
          24:
            level_vec_out = 64'b1111111111011110111111111101110111101111011111111111111001111111;
          25:
            level_vec_out = 64'b1111111111111110111111111101110111101111011111111111111001111111;
          26:
            level_vec_out = 64'b1111111111111110111111111101110111101111011111111111111101111111;
          27:
            level_vec_out = 64'b1111111111111110111111111101110111101111011111111111111101111111;
          28:
            level_vec_out = 64'b1111111111111111111111111101110111101111011111111111111101111111;
          29:
            level_vec_out = 64'b1111111111111111111111111111111111101111011111111111111101111111;
          30:
            level_vec_out = 64'b1111111111111111111111111111111111101111011111111111111101111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111101111011111111111111101111111;
        endcase
      1:
        case (frame_id)
          0:
            level_vec_out = 64'b0011110001000100101010000000010110101101010110011100110001101111;
          1:
            level_vec_out = 64'b0011110001001101101010010001010110101101010110011100110011101111;
          2:
            level_vec_out = 64'b0011110001001101101010010001010110101101110110011100110011101111;
          3:
            level_vec_out = 64'b0111110001001101101010010001010110101101110110011100110011101111;
          4:
            level_vec_out = 64'b0111110001001101101010010001010110101101110110011100110011101111;
          5:
            level_vec_out = 64'b0111110001001101101010010001110110101101110110011100110011101111;
          6:
            level_vec_out = 64'b0111110001001101101010110101110110101101110110011100110011101111;
          7:
            level_vec_out = 64'b0111110001001111101010110101110110101101111110011100110011101111;
          8:
            level_vec_out = 64'b0111110001001111101110110101110110101101111110011100110111101111;
          9:
            level_vec_out = 64'b0111110001001111101110110101110110101111111110011100110111101111;
          10:
            level_vec_out = 64'b0111110011001111101110110101110110101111111110011100110111101111;
          11:
            level_vec_out = 64'b0111110011001111101110110101110111101111111110011100110111101111;
          12:
            level_vec_out = 64'b0111110011001111101110110101110111101111111110011100110111101111;
          13:
            level_vec_out = 64'b0111110011001111101110110101111111101111111110111100110111101111;
          14:
            level_vec_out = 64'b0111110011001111101110110101111111101111111110111100110111101111;
          15:
            level_vec_out = 64'b0111110011001111111110110101111111101111111110111100111111101111;
          16:
            level_vec_out = 64'b0111110011001111111110110101111111101111111110111100111111101111;
          17:
            level_vec_out = 64'b0111111011011111111110110101111111101111111110111100111111101111;
          18:
            level_vec_out = 64'b0111111011011111111110110101111111101111111110111101111111101111;
          19:
            level_vec_out = 64'b0111111011011111111110110101111111101111111110111101111111111111;
          20:
            level_vec_out = 64'b0111111011011111111110110101111111101111111110111101111111111111;
          21:
            level_vec_out = 64'b0111111011011111111111110111111111101111111110111101111111111111;
          22:
            level_vec_out = 64'b0111111011011111111111110111111111101111111110111101111111111111;
          23:
            level_vec_out = 64'b1111111011011111111111110111111111101111111110111101111111111111;
          24:
            level_vec_out = 64'b1111111011011111111111110111111111111111111110111101111111111111;
          25:
            level_vec_out = 64'b1111111011011111111111110111111111111111111110111101111111111111;
          26:
            level_vec_out = 64'b1111111011011111111111110111111111111111111111111101111111111111;
          27:
            level_vec_out = 64'b1111111011011111111111110111111111111111111111111101111111111111;
          28:
            level_vec_out = 64'b1111111011011111111111110111111111111111111111111101111111111111;
          29:
            level_vec_out = 64'b1111111011011111111111110111111111111111111111111111111111111111;
          30:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        endcase
      2:
        case (frame_id)
          0:
            level_vec_out = 64'b1001010000000001011000110001100001100100000011111111101101000011;
          1:
            level_vec_out = 64'b1001010000000001011000110001110001100100000011111111101101000011;
          2:
            level_vec_out = 64'b1001010000000001011000110001110001100100000011111111101101000011;
          3:
            level_vec_out = 64'b1001010000000001011000110011110001100101000011111111101101000011;
          4:
            level_vec_out = 64'b1101010000000001011000110011110001100101000011111111101101000011;
          5:
            level_vec_out = 64'b1101010000000001011000110111110001100101000011111111101101001011;
          6:
            level_vec_out = 64'b1101010010000001011000110111110001100101000011111111101101001011;
          7:
            level_vec_out = 64'b1101010010000001011000110111110001100101000011111111101101001011;
          8:
            level_vec_out = 64'b1101010010000001011000110111110001100101000011111111101101001011;
          9:
            level_vec_out = 64'b1101010010010001011000110111110001100101000011111111101101001011;
          10:
            level_vec_out = 64'b1101010010010001011010110111110001100101000011111111101101001011;
          11:
            level_vec_out = 64'b1101010010110001011010110111110001100101000011111111101101001011;
          12:
            level_vec_out = 64'b1101010010110001011010110111110001100111000011111111101101001011;
          13:
            level_vec_out = 64'b1101010010110001011010110111110001100111000011111111101101001011;
          14:
            level_vec_out = 64'b1101010010110101011010110111110001100111000011111111101101011011;
          15:
            level_vec_out = 64'b1101010010110101011010110111110001100111000011111111101101011011;
          16:
            level_vec_out = 64'b1101010010110101011010110111110001101111000011111111101101011011;
          17:
            level_vec_out = 64'b1101010010110101011010110111110001101111000011111111111101011011;
          18:
            level_vec_out = 64'b1101010010110101011010110111110001101111000111111111111101111011;
          19:
            level_vec_out = 64'b1101010010110101011010110111110001101111000111111111111101111111;
          20:
            level_vec_out = 64'b1101011010110101011010110111110001111111010111111111111101111111;
          21:
            level_vec_out = 64'b1111011010110101011010110111111001111111010111111111111101111111;
          22:
            level_vec_out = 64'b1111011010110101011010110111111001111111010111111111111101111111;
          23:
            level_vec_out = 64'b1111011010110101011010110111111001111111010111111111111101111111;
          24:
            level_vec_out = 64'b1111011010110101011011110111111001111111010111111111111111111111;
          25:
            level_vec_out = 64'b1111111110110101011011110111111001111111010111111111111111111111;
          26:
            level_vec_out = 64'b1111111110110101011011110111111001111111010111111111111111111111;
          27:
            level_vec_out = 64'b1111111110110101011111110111111001111111110111111111111111111111;
          28:
            level_vec_out = 64'b1111111110110101011111110111111101111111110111111111111111111111;
          29:
            level_vec_out = 64'b1111111110110101011111110111111101111111110111111111111111111111;
          30:
            level_vec_out = 64'b1111111110110101011111110111111101111111110111111111111111111111;
          31:
            level_vec_out = 64'b1111111110111101111111110111111111111111111111111111111111111111;
        endcase
      3:
        case (frame_id)
          0:
            level_vec_out = 64'b0111000001100010100101001001100001011111000111100100010100010111;
          1:
            level_vec_out = 64'b0111000001100010100101001001101001011111000111100100010100010111;
          2:
            level_vec_out = 64'b0111000011100010100101001001101001011111000111100100010100010111;
          3:
            level_vec_out = 64'b0111000011100010100101001001101001011111000111100100010100010111;
          4:
            level_vec_out = 64'b0111000011100010100101001101101001011111010111100100010100010111;
          5:
            level_vec_out = 64'b0111000011100010100101001101101001011111010111100100010100010111;
          6:
            level_vec_out = 64'b0111000111100010100101001101101001011111010111100100010100010111;
          7:
            level_vec_out = 64'b0111000111100010100101001101101001011111010111100100010100010111;
          8:
            level_vec_out = 64'b0111000111100010100101001101101001011111011111110100010100010111;
          9:
            level_vec_out = 64'b0111000111100010110101001111101001011111011111110100010100010111;
          10:
            level_vec_out = 64'b0111000111100010110111001111101001011111011111110100010100010111;
          11:
            level_vec_out = 64'b0111000111100011110111001111101001011111011111110100010100011111;
          12:
            level_vec_out = 64'b0111000111100011110111001111101001011111011111110100010100011111;
          13:
            level_vec_out = 64'b0111000111100011110111001111101001011111011111110100010110011111;
          14:
            level_vec_out = 64'b0111000111100011110111001111101011011111111111110100010110011111;
          15:
            level_vec_out = 64'b0111001111100011110111001111101011011111111111110100010110011111;
          16:
            level_vec_out = 64'b1111101111100011110111001111101011011111111111110100010110011111;
          17:
            level_vec_out = 64'b1111101111100011110111001111101011011111111111110100010110011111;
          18:
            level_vec_out = 64'b1111101111100011110111101111101011011111111111110100010110011111;
          19:
            level_vec_out = 64'b1111101111100011110111101111101011011111111111110100010110011111;
          20:
            level_vec_out = 64'b1111101111100011110111101111101011011111111111110100010110011111;
          21:
            level_vec_out = 64'b1111111111100011110111111111101011111111111111110100010110011111;
          22:
            level_vec_out = 64'b1111111111100011110111111111101011111111111111110100011110011111;
          23:
            level_vec_out = 64'b1111111111110011110111111111101011111111111111110100011110011111;
          24:
            level_vec_out = 64'b1111111111110011111111111111101011111111111111110101011110011111;
          25:
            level_vec_out = 64'b1111111111111011111111111111111011111111111111110101011111011111;
          26:
            level_vec_out = 64'b1111111111111011111111111111111011111111111111110101011111011111;
          27:
            level_vec_out = 64'b1111111111111011111111111111111011111111111111111101011111011111;
          28:
            level_vec_out = 64'b1111111111111011111111111111111011111111111111111101011111011111;
          29:
            level_vec_out = 64'b1111111111111011111111111111111111111111111111111101011111111111;
          30:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111101011111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        endcase
      4:
        case (frame_id)
          0:
            level_vec_out = 64'b0001101100011100001101111011010110001001001000010101111011101100;
          1:
            level_vec_out = 64'b0001101100011100001101111011010110001001001000010101111011101100;
          2:
            level_vec_out = 64'b0001101100011100001101111011010110001001001000010101111011101100;
          3:
            level_vec_out = 64'b0001111100011100001101111011011110001001001000010101111011101100;
          4:
            level_vec_out = 64'b0001111100011100001101111011111110001001001000010101111011101101;
          5:
            level_vec_out = 64'b0001111100011100001101111011111110001001001000010101111011101101;
          6:
            level_vec_out = 64'b0001111100011101001101111011111110001001001010010101111011101101;
          7:
            level_vec_out = 64'b0001111100011101001101111011111110001001011010010101111111101101;
          8:
            level_vec_out = 64'b0001111100011101001101111011111110001001011010011101111111101101;
          9:
            level_vec_out = 64'b0111111100011101001101111011111110001001011010011101111111101101;
          10:
            level_vec_out = 64'b0111111100011101001101111011111110101001011010011101111111111101;
          11:
            level_vec_out = 64'b0111111100011101001101111011111110101001011010011101111111111101;
          12:
            level_vec_out = 64'b0111111100011111101101111111111110101001011010011101111111111101;
          13:
            level_vec_out = 64'b0111111110011111101111111111111110101001111010011101111111111101;
          14:
            level_vec_out = 64'b0111111110011111101111111111111110101001111010011111111111111101;
          15:
            level_vec_out = 64'b0111111110011111101111111111111110101001111010011111111111111101;
          16:
            level_vec_out = 64'b0111111110011111101111111111111110101001111010011111111111111101;
          17:
            level_vec_out = 64'b0111111110011111101111111111111110101001111110011111111111111101;
          18:
            level_vec_out = 64'b0111111110011111101111111111111110101001111110011111111111111101;
          19:
            level_vec_out = 64'b0111111110011111111111111111111110101001111110011111111111111101;
          20:
            level_vec_out = 64'b0111111110011111111111111111111110101101111110011111111111111101;
          21:
            level_vec_out = 64'b0111111110011111111111111111111110101101111110011111111111111101;
          22:
            level_vec_out = 64'b0111111110011111111111111111111111101101111110011111111111111101;
          23:
            level_vec_out = 64'b0111111110011111111111111111111111101101111110011111111111111101;
          24:
            level_vec_out = 64'b0111111110011111111111111111111111111101111110011111111111111111;
          25:
            level_vec_out = 64'b0111111110011111111111111111111111111101111110011111111111111111;
          26:
            level_vec_out = 64'b0111111110011111111111111111111111111101111110111111111111111111;
          27:
            level_vec_out = 64'b0111111110011111111111111111111111111111111110111111111111111111;
          28:
            level_vec_out = 64'b1111111111011111111111111111111111111111111110111111111111111111;
          29:
            level_vec_out = 64'b1111111111011111111111111111111111111111111110111111111111111111;
          30:
            level_vec_out = 64'b1111111111011111111111111111111111111111111110111111111111111111;
          31:
            level_vec_out = 64'b1111111111011111111111111111111111111111111111111111111111111111;
        endcase
      5:
        case (frame_id)
          0:
            level_vec_out = 64'b0000011001001000001010011110010111101111101000100010100110010111;
          1:
            level_vec_out = 64'b0000011001001000001010011110010111101111101000100010110110010111;
          2:
            level_vec_out = 64'b0000011001001000001010011110010111101111101000100010110110010111;
          3:
            level_vec_out = 64'b0000011001001000001010011110010111101111101000100110110110010111;
          4:
            level_vec_out = 64'b0000011001001000001010011110010111101111101000100111110110010111;
          5:
            level_vec_out = 64'b0000111001001000001010011110010111101111101000100111110110010111;
          6:
            level_vec_out = 64'b0000111001001000001010011110010111101111101000100111110110010111;
          7:
            level_vec_out = 64'b0000111001001000101010011110010111101111101000100111110110010111;
          8:
            level_vec_out = 64'b0000111001001000101010011110010111101111101000100111110111011111;
          9:
            level_vec_out = 64'b0000111001001000101010011110010111101111101000100111110111011111;
          10:
            level_vec_out = 64'b0000111001001100101010011110010111101111101000100111110111011111;
          11:
            level_vec_out = 64'b0000111001001100101010011110010111101111101001100111110111011111;
          12:
            level_vec_out = 64'b0001111001001100101010011110011111101111101001100111110111011111;
          13:
            level_vec_out = 64'b0001111001001100101010011110011111101111101001100111110111011111;
          14:
            level_vec_out = 64'b0001111001001100101010011110011111101111101101100111110111011111;
          15:
            level_vec_out = 64'b0001111101001100101010011110111111101111101101110111110111011111;
          16:
            level_vec_out = 64'b0001111101011100101010011110111111101111101111110111110111011111;
          17:
            level_vec_out = 64'b0001111101011100111011011110111111101111101111110111110111011111;
          18:
            level_vec_out = 64'b0001111111011100111011011110111111101111101111110111110111011111;
          19:
            level_vec_out = 64'b0101111111011101111011011110111111101111101111110111110111011111;
          20:
            level_vec_out = 64'b0111111111011101111011011110111111101111101111110111110111011111;
          21:
            level_vec_out = 64'b0111111111011101111011011110111111101111101111110111110111011111;
          22:
            level_vec_out = 64'b0111111111111111111011011110111111101111101111110111111111011111;
          23:
            level_vec_out = 64'b0111111111111111111011011110111111101111111111110111111111011111;
          24:
            level_vec_out = 64'b0111111111111111111011011110111111101111111111110111111111011111;
          25:
            level_vec_out = 64'b0111111111111111111011011110111111101111111111110111111111011111;
          26:
            level_vec_out = 64'b1111111111111111111011111110111111101111111111110111111111011111;
          27:
            level_vec_out = 64'b1111111111111111111011111110111111101111111111110111111111011111;
          28:
            level_vec_out = 64'b1111111111111111111011111111111111111111111111110111111111011111;
          29:
            level_vec_out = 64'b1111111111111111111011111111111111111111111111111111111111111111;
          30:
            level_vec_out = 64'b1111111111111111111011111111111111111111111111111111111111111111;
          31:
            level_vec_out = 64'b1111111111111111111011111111111111111111111111111111111111111111;
        endcase
      6:
        case (frame_id)
          0:
            level_vec_out = 64'b1111011111001010001111011111010000011111111001101100011111011000;
          1:
            level_vec_out = 64'b1111011111001010001111011111010000011111111001101100011111011000;
          2:
            level_vec_out = 64'b1111011111001011001111011111010000011111111001101100011111011101;
          3:
            level_vec_out = 64'b1111011111001011001111011111010000011111111001101100011111011101;
          4:
            level_vec_out = 64'b1111011111001011001111011111010000011111111001101100011111011101;
          5:
            level_vec_out = 64'b1111011111001111001111011111010000011111111001101100011111011101;
          6:
            level_vec_out = 64'b1111011111001111001111011111010100011111111001111100011111011101;
          7:
            level_vec_out = 64'b1111011111001111001111011111010100011111111001111100011111011101;
          8:
            level_vec_out = 64'b1111011111001111001111011111010100011111111001111100111111011101;
          9:
            level_vec_out = 64'b1111011111001111001111011111010100011111111001111110111111011101;
          10:
            level_vec_out = 64'b1111011111001111001111011111010100011111111001111110111111011101;
          11:
            level_vec_out = 64'b1111011111001111101111011111010100011111111001111110111111011101;
          12:
            level_vec_out = 64'b1111011111001111101111011111010100011111111001111110111111011101;
          13:
            level_vec_out = 64'b1111011111001111101111011111010100011111111001111110111111011101;
          14:
            level_vec_out = 64'b1111011111001111101111011111010100011111111001111110111111011101;
          15:
            level_vec_out = 64'b1111011111001111101111011111010100011111111001111110111111011101;
          16:
            level_vec_out = 64'b1111011111011111101111011111010100011111111001111110111111011101;
          17:
            level_vec_out = 64'b1111011111011111101111011111010100011111111001111110111111011101;
          18:
            level_vec_out = 64'b1111011111011111101111011111010100111111111001111110111111011101;
          19:
            level_vec_out = 64'b1111011111011111101111011111010100111111111011111110111111011111;
          20:
            level_vec_out = 64'b1111011111011111101111011111010100111111111011111110111111011111;
          21:
            level_vec_out = 64'b1111011111011111101111011111010100111111111011111111111111011111;
          22:
            level_vec_out = 64'b1111111111011111101111011111010100111111111011111111111111011111;
          23:
            level_vec_out = 64'b1111111111011111101111011111110100111111111011111111111111011111;
          24:
            level_vec_out = 64'b1111111111011111101111011111110100111111111011111111111111011111;
          25:
            level_vec_out = 64'b1111111111011111101111011111110100111111111011111111111111011111;
          26:
            level_vec_out = 64'b1111111111111111101111011111110101111111111011111111111111011111;
          27:
            level_vec_out = 64'b1111111111111111111111011111110101111111111111111111111111011111;
          28:
            level_vec_out = 64'b1111111111111111111111111111110101111111111111111111111111011111;
          29:
            level_vec_out = 64'b1111111111111111111111111111110101111111111111111111111111111111;
          30:
            level_vec_out = 64'b1111111111111111111111111111110111111111111111111111111111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        endcase
      7:
        case (frame_id)
          0:
            level_vec_out = 64'b1111011010111000110110000010101010011111001110001011001000111010;
          1:
            level_vec_out = 64'b1111011010111000110110000010101010011111001110001011001000111010;
          2:
            level_vec_out = 64'b1111011010111000110110000010101010011111001110001011001000111010;
          3:
            level_vec_out = 64'b1111011010111000110110000010101010011111001110001011001000111010;
          4:
            level_vec_out = 64'b1111011010111000110110000110101010011111001110001011001001111010;
          5:
            level_vec_out = 64'b1111011010111000110110000110101110011111001110101011001001111010;
          6:
            level_vec_out = 64'b1111011010111000110110000110101110011111001110101011001001111010;
          7:
            level_vec_out = 64'b1111011010111000110110000110101110011111001110101011001001111010;
          8:
            level_vec_out = 64'b1111011010111000110110000110101110011111001110101011001001111010;
          9:
            level_vec_out = 64'b1111011010111000110110000110101110011111001110101011001001111010;
          10:
            level_vec_out = 64'b1111011010111000110110010110101110011111001111101011001001111010;
          11:
            level_vec_out = 64'b1111011010111000110110010110101110011111001111101011001001111010;
          12:
            level_vec_out = 64'b1111011010111000110110010110101110011111001111101011001001111110;
          13:
            level_vec_out = 64'b1111011010111000110110010110101110011111001111101011011001111110;
          14:
            level_vec_out = 64'b1111011010111000110111010110101110011111001111111011011001111110;
          15:
            level_vec_out = 64'b1111011010111000110111010110101110011111001111111011011001111110;
          16:
            level_vec_out = 64'b1111011010111000110111010110101110111111001111111011011001111110;
          17:
            level_vec_out = 64'b1111011110111000110111010110101110111111001111111011011001111110;
          18:
            level_vec_out = 64'b1111011110111000110111010110101110111111001111111111011001111110;
          19:
            level_vec_out = 64'b1111011110111000110111010110101110111111101111111111011001111110;
          20:
            level_vec_out = 64'b1111011110111100110111011110101110111111101111111111011001111110;
          21:
            level_vec_out = 64'b1111011110111100110111011110101110111111101111111111011001111110;
          22:
            level_vec_out = 64'b1111011110111100110111011110101111111111101111111111011001111110;
          23:
            level_vec_out = 64'b1111011110111111110111111110101111111111101111111111011001111110;
          24:
            level_vec_out = 64'b1111011110111111110111111110101111111111101111111111011001111111;
          25:
            level_vec_out = 64'b1111011111111111110111111110101111111111101111111111011101111111;
          26:
            level_vec_out = 64'b1111011111111111111111111110101111111111101111111111011101111111;
          27:
            level_vec_out = 64'b1111111111111111111111111110101111111111111111111111011101111111;
          28:
            level_vec_out = 64'b1111111111111111111111111110111111111111111111111111011101111111;
          29:
            level_vec_out = 64'b1111111111111111111111111110111111111111111111111111011101111111;
          30:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        endcase
    endcase
  end
endmodule