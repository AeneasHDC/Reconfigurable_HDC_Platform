----
 -- @file level_hvec_gen_hdl.hpp
 -- @brief This script generates HDL code for generating high-dimensional LEVEL vectors.
 -- It is a novel method; for more information, please refer to our paper.
 --
 -- @author Saeid Jamili and Marco Angioli
 -- @note Author names are listed in alphabetical order.
 -- @email <saeid.jamili@uniroma1.it>
 -- @email <marco.angioli@uniroma1.it>
 --
 -- @contributors
 --
 -- @date Created: 24th July 2023
 -- @date Last Updated: 23th August 2023
 --
 -- @version 1.0.0
 --
 -- @institute Sapienza University of Rome
 -- @cite https://doi.org/10.xxxx/yyyyy
 --
 -- @section DEPENDENCIES
 -- - Dependency1: Description or version details.
 -- - Dependency2: Description or version details.
 --
 -- @section LICENSE
 -- This file is part of the Aeneas HyperCompute Platform.
 --
 -- Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 --
 -- @section CHANGELOG
 -- @version 1.0.0-dev - 23th August 2023
 -- - Initial release
 --
 -- @todo
 -- - Complete level vector generator function
 -- - Add training
 --
 -- @see
 -- -
 -- -
 -- -
 --
 --

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity level_vec_gen is
    Port ( level_vec_out : out  STD_LOGIC_VECTOR (63 downto 0);
           frame_index : in  STD_LOGIC_VECTOR (2 downto 0);
           frame_id : in  STD_LOGIC_VECTOR (4 downto 0));
end level_vec_gen;

architecture Behavioral of level_vec_gen is
begin
    process (frame_index, frame_id)
    begin
        -- Update this function to match your requirements
        case frame_index is
            when "000" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1111110101000000111110100100110111110100110000111000110010000011";
                    when "00001" => level_vec_out <= "1111110101000000111110100100110111110100110000111000110010000011";
                    when "00010" => level_vec_out <= "1111110101000100111110100110110111110100110000111000110010000011";
                    when "00011" => level_vec_out <= "1111110101010100111110100110110111111100110000111000110010000011";
                    when "00100" => level_vec_out <= "1111110101010100111110100110110111111100110000111001110010010011";
                    when "00101" => level_vec_out <= "1111110101010101111110100110110111111100110000111001110010010011";
                    when "00110" => level_vec_out <= "1111110101010101111110100110110111111100110000111001111010010011";
                    when "00111" => level_vec_out <= "1111110101110101111110100110110111111100110000111001111010010011";
                    when "01000" => level_vec_out <= "1111110101110101111110100110110111111100110000111001111010010111";
                    when "01001" => level_vec_out <= "1111110101110101111110100110110111111100110000111001111010010111";
                    when "01010" => level_vec_out <= "1111110101110101111110100110110111111100110000111001111010010111";
                    when "01011" => level_vec_out <= "1111110101110101111110100110110111111100110000111001111110011111";
                    when "01100" => level_vec_out <= "1111110101111101111110100110110111111100110000111001111110011111";
                    when "01101" => level_vec_out <= "1111110101111101111110100110110111111100110000111001111110011111";
                    when "01110" => level_vec_out <= "1111110101111101111110100110110111111101110010111001111110011111";
                    when "01111" => level_vec_out <= "1111110101111101111110110110110111111101110010111001111110011111";
                    when "10000" => level_vec_out <= "1111110101111101111110110110110111111111110010111001111110011111";
                    when "10001" => level_vec_out <= "1111110101111101111110111110110111111111110010111001111110011111";
                    when "10010" => level_vec_out <= "1111111101111101111110111110110111111111110010111101111110011111";
                    when "10011" => level_vec_out <= "1111111101111101111110111110110111111111110010111101111110111111";
                    when "10100" => level_vec_out <= "1111111101111101111110111110110111111111110010111101111110111111";
                    when "10101" => level_vec_out <= "1111111101111101111110111110110111111111110010111101111110111111";
                    when "10110" => level_vec_out <= "1111111101111101111110111110110111111111110011111101111110111111";
                    when "10111" => level_vec_out <= "1111111101111111111110111110110111111111110011111101111110111111";
                    when "11000" => level_vec_out <= "1111111101111111111110111110110111111111111011111101111110111111";
                    when "11001" => level_vec_out <= "1111111111111111111111111110110111111111111011111101111110111111";
                    when "11010" => level_vec_out <= "1111111111111111111111111110110111111111111011111101111110111111";
                    when "11011" => level_vec_out <= "1111111111111111111111111110110111111111111011111101111111111111";
                    when "11100" => level_vec_out <= "1111111111111111111111111110111111111111111011111101111111111111";
                    when "11101" => level_vec_out <= "1111111111111111111111111110111111111111111011111101111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111111011111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111011111111111111111111";
                when others => null;
                end case;
            when "001" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0111001001101101110000011010100100010001111110000100100011011010";
                    when "00001" => level_vec_out <= "0111001001101101110100011010101100010001111110000100100011011010";
                    when "00010" => level_vec_out <= "0111001001101101110100011010101100010001111110000100100011011011";
                    when "00011" => level_vec_out <= "0111001001101101110100011010101100010001111110000100100011011011";
                    when "00100" => level_vec_out <= "0111001001101101110100011010101100010001111110000100100011011011";
                    when "00101" => level_vec_out <= "0111001001101101110100011010101100011001111110000100100011111011";
                    when "00110" => level_vec_out <= "0111001001101101110100011010101100011001111110000100100011111011";
                    when "00111" => level_vec_out <= "0111001001101101110100011010101100011001111110000100100011111011";
                    when "01000" => level_vec_out <= "0111101001101101110100011010101100011001111110000100111011111011";
                    when "01001" => level_vec_out <= "0111101001101101110100011010101100011001111110000100111011111011";
                    when "01010" => level_vec_out <= "0111101001101111110100011111101100011001111110000100111011111011";
                    when "01011" => level_vec_out <= "0111101001101111110100011111101100011001111110000100111011111011";
                    when "01100" => level_vec_out <= "0111101001101111110100011111101110011001111110000100111011111011";
                    when "01101" => level_vec_out <= "0111101001101111111100011111101110011001111110110100111011111011";
                    when "01110" => level_vec_out <= "0111111001101111111100011111101110011001111111110100111011111011";
                    when "01111" => level_vec_out <= "0111111001101111111100011111101110011001111111110100111011111011";
                    when "10000" => level_vec_out <= "0111111001101111111100011111101110011001111111110110111011111011";
                    when "10001" => level_vec_out <= "0111111001101111111100011111101110011001111111110110111011111011";
                    when "10010" => level_vec_out <= "0111111001101111111100011111101110011001111111110110111011111111";
                    when "10011" => level_vec_out <= "0111111001101111111100011111101110011011111111110110111011111111";
                    when "10100" => level_vec_out <= "0111111001101111111100011111101111011011111111110111111011111111";
                    when "10101" => level_vec_out <= "0111111101101111111100011111101111011111111111110111111011111111";
                    when "10110" => level_vec_out <= "0111111101101111111100011111101111011111111111110111111011111111";
                    when "10111" => level_vec_out <= "0111111111101111111100011111101111011111111111110111111011111111";
                    when "11000" => level_vec_out <= "0111111111101111111100011111101111011111111111111111111011111111";
                    when "11001" => level_vec_out <= "0111111111101111111110011111101111011111111111111111111011111111";
                    when "11010" => level_vec_out <= "0111111111101111111110011111111111011111111111111111111011111111";
                    when "11011" => level_vec_out <= "0111111111101111111111011111111111011111111111111111111011111111";
                    when "11100" => level_vec_out <= "0111111111101111111111011111111111011111111111111111111011111111";
                    when "11101" => level_vec_out <= "0111111111101111111111111111111111011111111111111111111011111111";
                    when "11110" => level_vec_out <= "0111111111111111111111111111111111111111111111111111111011111111";
                    when "11111" => level_vec_out <= "0111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "010" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0011111000111100011010100100011110101110110100001000000100001000";
                    when "00001" => level_vec_out <= "0011111000111100011010100100011110101110110100001000000100001100";
                    when "00010" => level_vec_out <= "1011111000111100011010100100011110101110110100001000000100001101";
                    when "00011" => level_vec_out <= "1011111000111100011010100100011110101110110100001001000100001101";
                    when "00100" => level_vec_out <= "1011111000111100011010100100011110101110110100001001000100001101";
                    when "00101" => level_vec_out <= "1011111000111110011010100100011110101110110100001001000100101101";
                    when "00110" => level_vec_out <= "1011111001111110011010100100011110101110110100001001000100101101";
                    when "00111" => level_vec_out <= "1011111001111110011010100100011110101110110100001001000100101111";
                    when "01000" => level_vec_out <= "1011111001111110011010101100011110101110110100001001000100101111";
                    when "01001" => level_vec_out <= "1011111001111110011010101100011110101110110100001001000100101111";
                    when "01010" => level_vec_out <= "1011111001111110011010101100011110101110110100001101000100111111";
                    when "01011" => level_vec_out <= "1011111001111110011010101100011110101110110100001101000100111111";
                    when "01100" => level_vec_out <= "1011111001111110011010101100011110101110110110001101000100111111";
                    when "01101" => level_vec_out <= "1011111001111110011010111100011110101110110111001101000100111111";
                    when "01110" => level_vec_out <= "1011111001111110011010111100111110101111110111001101000100111111";
                    when "01111" => level_vec_out <= "1011111001111110011010111100111110101111110111001101000101111111";
                    when "10000" => level_vec_out <= "1011111001111110011011111100111110111111110111001101000101111111";
                    when "10001" => level_vec_out <= "1011111011111110011011111101111110111111110111001101000101111111";
                    when "10010" => level_vec_out <= "1011111011111110011011111101111110111111110111011101000101111111";
                    when "10011" => level_vec_out <= "1011111111111110011011111101111111111111110111011101000101111111";
                    when "10100" => level_vec_out <= "1011111111111110011011111101111111111111110111011101000101111111";
                    when "10101" => level_vec_out <= "1011111111111110011011111101111111111111110111111101100101111111";
                    when "10110" => level_vec_out <= "1011111111111110011111111101111111111111110111111101110101111111";
                    when "10111" => level_vec_out <= "1011111111111110011111111101111111111111110111111101110101111111";
                    when "11000" => level_vec_out <= "1011111111111110111111111101111111111111110111111101110101111111";
                    when "11001" => level_vec_out <= "1011111111111110111111111101111111111111110111111101110101111111";
                    when "11010" => level_vec_out <= "1011111111111110111111111101111111111111110111111101110101111111";
                    when "11011" => level_vec_out <= "1011111111111110111111111101111111111111110111111101110101111111";
                    when "11100" => level_vec_out <= "1011111111111110111111111101111111111111111111111101111111111111";
                    when "11101" => level_vec_out <= "1011111111111110111111111111111111111111111111111101111111111111";
                    when "11110" => level_vec_out <= "1011111111111111111111111111111111111111111111111101111111111111";
                    when "11111" => level_vec_out <= "1011111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "011" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1101010011010000000100111001111001011111100010111101001110111111";
                    when "00001" => level_vec_out <= "1101010011010000000100111001111001011111100010111101001110111111";
                    when "00010" => level_vec_out <= "1101010011010000000110111001111001011111100010111101001110111111";
                    when "00011" => level_vec_out <= "1101010011010000000110111001111001011111100110111101001110111111";
                    when "00100" => level_vec_out <= "1101010011010000010110111001111001011111100110111101001110111111";
                    when "00101" => level_vec_out <= "1101010011010000010110111001111001011111100110111101001110111111";
                    when "00110" => level_vec_out <= "1101010011010100010110111001111001011111100110111101001110111111";
                    when "00111" => level_vec_out <= "1101010011010100010110111101111001111111100110111101101110111111";
                    when "01000" => level_vec_out <= "1101010011010100010110111101111001111111100110111101101110111111";
                    when "01001" => level_vec_out <= "1101110011010100010110111101111001111111100110111101101110111111";
                    when "01010" => level_vec_out <= "1101110011010100010110111101111001111111100110111101101110111111";
                    when "01011" => level_vec_out <= "1101110011010100110110111101111001111111100110111111101110111111";
                    when "01100" => level_vec_out <= "1101110011010100110110111101111001111111100110111111101110111111";
                    when "01101" => level_vec_out <= "1101110011010100110110111101111001111111100110111111101110111111";
                    when "01110" => level_vec_out <= "1101110111010100110110111101111001111111100110111111101110111111";
                    when "01111" => level_vec_out <= "1101110111010100110110111101111001111111100110111111101110111111";
                    when "10000" => level_vec_out <= "1101110111010100110110111101111001111111100110111111101110111111";
                    when "10001" => level_vec_out <= "1101110111010100110110111101111001111111100110111111101110111111";
                    when "10010" => level_vec_out <= "1101110111010100110110111101111001111111100110111111101110111111";
                    when "10011" => level_vec_out <= "1101110111010100110110111101111001111111110110111111101110111111";
                    when "10100" => level_vec_out <= "1101111111010100111110111101111001111111110110111111101110111111";
                    when "10101" => level_vec_out <= "1101111111010100111110111101111001111111110110111111101110111111";
                    when "10110" => level_vec_out <= "1101111111010100111111111101111001111111110110111111101111111111";
                    when "10111" => level_vec_out <= "1101111111010100111111111101111001111111110110111111111111111111";
                    when "11000" => level_vec_out <= "1111111111010100111111111101111101111111110110111111111111111111";
                    when "11001" => level_vec_out <= "1111111111010110111111111101111101111111111110111111111111111111";
                    when "11010" => level_vec_out <= "1111111111010110111111111111111111111111111110111111111111111111";
                    when "11011" => level_vec_out <= "1111111111010111111111111111111111111111111110111111111111111111";
                    when "11100" => level_vec_out <= "1111111111010111111111111111111111111111111110111111111111111111";
                    when "11101" => level_vec_out <= "1111111111111111111111111111111111111111111110111111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when "100" =>
                case frame_id is
                    when "00000" => level_vec_out <= "1100011001101101000010101110011001011001101100110110111011010001";
                    when "00001" => level_vec_out <= "1100011001101101000010101110011001011001101100110111111011010001";
                    when "00010" => level_vec_out <= "1100011001101101000010101110011001011001101100110111111011010001";
                    when "00011" => level_vec_out <= "1100011001101101000010101110011101011001101100110111111011010001";
                    when "00100" => level_vec_out <= "1100011001101101000010101110011111011001101100110111111011010001";
                    when "00101" => level_vec_out <= "1100111001101101000010101110011111011001101100110111111011010001";
                    when "00110" => level_vec_out <= "1100111001101101000010101110011111011001101100110111111011010001";
                    when "00111" => level_vec_out <= "1100111001101101000010101110011111011001101100110111111011010101";
                    when "01000" => level_vec_out <= "1100111001101101001010101110011111011001101100110111111011010101";
                    when "01001" => level_vec_out <= "1100111111101101001010101110011111011001101110110111111011010101";
                    when "01010" => level_vec_out <= "1100111111101101001010101110011111011001101110110111111111010101";
                    when "01011" => level_vec_out <= "1100111111101101001010101110011111011001101110110111111111010101";
                    when "01100" => level_vec_out <= "1100111111101101001010101110011111011001101110110111111111010101";
                    when "01101" => level_vec_out <= "1110111111101101001010101110011111011001101110110111111111010101";
                    when "01110" => level_vec_out <= "1110111111101101001010101110011111011001101110110111111111010101";
                    when "01111" => level_vec_out <= "1110111111101111011010101110011111011001101110110111111111010101";
                    when "10000" => level_vec_out <= "1110111111101111011010101110011111011011101110110111111111010101";
                    when "10001" => level_vec_out <= "1110111111101111011010111110011111011011101110110111111111010101";
                    when "10010" => level_vec_out <= "1110111111101111011010111110011111011011101110110111111111010111";
                    when "10011" => level_vec_out <= "1110111111101111011010111110011111011011101110110111111111011111";
                    when "10100" => level_vec_out <= "1110111111101111011010111110011111111011101110110111111111011111";
                    when "10101" => level_vec_out <= "1110111111101111011010111110011111111011101110110111111111011111";
                    when "10110" => level_vec_out <= "1110111111101111011010111111011111111011101111110111111111011111";
                    when "10111" => level_vec_out <= "1110111111101111011011111111011111111011101111110111111111011111";
                    when "11000" => level_vec_out <= "1110111111101111011011111111011111111011101111110111111111011111";
                    when "11001" => level_vec_out <= "1110111111101111011011111111011111111011101111110111111111011111";
                    when "11010" => level_vec_out <= "1110111111101111011011111111111111111011111111110111111111011111";
                    when "11011" => level_vec_out <= "1110111111101111011011111111111111111111111111110111111111011111";
                    when "11100" => level_vec_out <= "1110111111111111011011111111111111111111111111110111111111011111";
                    when "11101" => level_vec_out <= "1110111111111111011011111111111111111111111111110111111111011111";
                    when "11110" => level_vec_out <= "1110111111111111111011111111111111111111111111111111111111011111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111111111111111111111111111111011111";
                when others => null;
                end case;
            when "101" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0011011111001000100101000000010011011110100001101010100100011100";
                    when "00001" => level_vec_out <= "0011011111001000100101000000010011011110100101101010100100011100";
                    when "00010" => level_vec_out <= "0011011111001000100101000000010011011110100101101010110100011100";
                    when "00011" => level_vec_out <= "0011011111001000100101000000010011011110100101101010110100011100";
                    when "00100" => level_vec_out <= "0011011111001000100101000000010011011110100101101110110100011100";
                    when "00101" => level_vec_out <= "0011011111001000100101000000010011011110100101101110110100011100";
                    when "00110" => level_vec_out <= "0011011111001000100101000000010011011110100101101110110100011100";
                    when "00111" => level_vec_out <= "0011011111001000100101000000010011111110100101101110110100011100";
                    when "01000" => level_vec_out <= "0011011111001000100101000000010011111110100101101110110100011100";
                    when "01001" => level_vec_out <= "0011011111001000100101000000010011111110100101101110110100011100";
                    when "01010" => level_vec_out <= "0011011111001000100101001000010011111110100101101110110100011100";
                    when "01011" => level_vec_out <= "0011011111001000100101001000011011111110100101101110111100011100";
                    when "01100" => level_vec_out <= "0011011111001000101101001100011011111110100101101110111100011100";
                    when "01101" => level_vec_out <= "0011011111001000101101001100011011111110100101101110111100011100";
                    when "01110" => level_vec_out <= "0011011111001000101101011100011011111110100101101110111100011100";
                    when "01111" => level_vec_out <= "0011111111001000101101011100111011111110100101101110111100111100";
                    when "10000" => level_vec_out <= "0011111111001001101101011100111011111110100101101110111100111100";
                    when "10001" => level_vec_out <= "0011111111001001101101011110111011111110100101101110111100111101";
                    when "10010" => level_vec_out <= "0011111111101001101101011110111011111110110101101110111110111101";
                    when "10011" => level_vec_out <= "0011111111101001101101011110111011111110110101101110111110111101";
                    when "10100" => level_vec_out <= "0011111111101001111101011110111111111110110101101110111110111101";
                    when "10101" => level_vec_out <= "0011111111111001111111111110111111111110110101101110111110111101";
                    when "10110" => level_vec_out <= "0011111111111001111111111110111111111110110101101110111110111111";
                    when "10111" => level_vec_out <= "0011111111111001111111111110111111111110110101101110111110111111";
                    when "11000" => level_vec_out <= "0011111111111011111111111110111111111110110101101110111111111111";
                    when "11001" => level_vec_out <= "0011111111111011111111111110111111111111110111101110111111111111";
                    when "11010" => level_vec_out <= "0011111111111011111111111111111111111111110111101110111111111111";
                    when "11011" => level_vec_out <= "1011111111111011111111111111111111111111110111101111111111111111";
                    when "11100" => level_vec_out <= "1011111111111011111111111111111111111111110111101111111111111111";
                    when "11101" => level_vec_out <= "1011111111111011111111111111111111111111110111101111111111111111";
                    when "11110" => level_vec_out <= "1011111111111011111111111111111111111111110111101111111111111111";
                    when "11111" => level_vec_out <= "1111111111111011111111111111111111111111111111101111111111111111";
                when others => null;
                end case;
            when "110" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0101111100101101000111010101111010001111101000001010000011100100";
                    when "00001" => level_vec_out <= "0101111100101101000111010101111010011111101000001110000011100100";
                    when "00010" => level_vec_out <= "0101111100101101000111010101111010011111101000001110000011100100";
                    when "00011" => level_vec_out <= "0101111100101101000111010101111010011111101000001110000011100100";
                    when "00100" => level_vec_out <= "0111111100101101000111010101111011011111101000001110000011100100";
                    when "00101" => level_vec_out <= "0111111100101101000111011101111011011111101000001110000011100100";
                    when "00110" => level_vec_out <= "0111111100101101000111011101111011011111101000001110100111100110";
                    when "00111" => level_vec_out <= "0111111100101101000111011101111011011111101000001110100111100110";
                    when "01000" => level_vec_out <= "0111111100101101000111011101111011011111101000001110100111100110";
                    when "01001" => level_vec_out <= "0111111111101101000111011101111011011111101010001110100111100110";
                    when "01010" => level_vec_out <= "0111111111101101000111011101111011011111101010001110100111110110";
                    when "01011" => level_vec_out <= "0111111111101101000111011101111011011111101010001110100111111110";
                    when "01100" => level_vec_out <= "0111111111101101000111011111111011011111111010001110100111111110";
                    when "01101" => level_vec_out <= "0111111111101101000111011111111011011111111011001110100111111110";
                    when "01110" => level_vec_out <= "0111111111101101000111011111111011011111111011001110100111111110";
                    when "01111" => level_vec_out <= "0111111111101101000111011111111011011111111011001110100111111110";
                    when "10000" => level_vec_out <= "0111111111101101000111011111111011011111111011001110100111111111";
                    when "10001" => level_vec_out <= "0111111111101101011111011111111011011111111011001110100111111111";
                    when "10010" => level_vec_out <= "0111111111101101011111011111111011011111111011001110100111111111";
                    when "10011" => level_vec_out <= "1111111111101101011111111111111011011111111011001110100111111111";
                    when "10100" => level_vec_out <= "1111111111101101011111111111111011011111111011001110100111111111";
                    when "10101" => level_vec_out <= "1111111111101101011111111111111011011111111011001110100111111111";
                    when "10110" => level_vec_out <= "1111111111101101011111111111111011011111111011001110100111111111";
                    when "10111" => level_vec_out <= "1111111111101101011111111111111011011111111011001110100111111111";
                    when "11000" => level_vec_out <= "1111111111101101011111111111111011011111111111001110100111111111";
                    when "11001" => level_vec_out <= "1111111111101101011111111111111011011111111111001110100111111111";
                    when "11010" => level_vec_out <= "1111111111101101011111111111111011111111111111001110100111111111";
                    when "11011" => level_vec_out <= "1111111111101101011111111111111011111111111111111110100111111111";
                    when "11100" => level_vec_out <= "1111111111111101011111111111111011111111111111111110100111111111";
                    when "11101" => level_vec_out <= "1111111111111111111111111111111011111111111111111110101111111111";
                    when "11110" => level_vec_out <= "1111111111111111111111111111111011111111111111111110101111111111";
                    when "11111" => level_vec_out <= "1111111111111111111111111111111011111111111111111111111111111111";
                when others => null;
                end case;
            when "111" =>
                case frame_id is
                    when "00000" => level_vec_out <= "0011011011100110111011100000010101111001111000010010100111010110";
                    when "00001" => level_vec_out <= "0011011011100110111011100010010101111001111000010010100111010110";
                    when "00010" => level_vec_out <= "0011011011100110111011100010010101111001111000010010101111010110";
                    when "00011" => level_vec_out <= "0011011011101110111011100010010101111101111000110010101111010110";
                    when "00100" => level_vec_out <= "0011011011101110111011100010010101111101111001110010101111010110";
                    when "00101" => level_vec_out <= "0011011011101110111011100010010101111101111001111010101111010110";
                    when "00110" => level_vec_out <= "0111011011101111111011100010010101111101111001111010101111010110";
                    when "00111" => level_vec_out <= "0111111011101111111011100010010101111101111001111010101111010110";
                    when "01000" => level_vec_out <= "0111111111111111111011100010010101111101111001111010101111010110";
                    when "01001" => level_vec_out <= "0111111111111111111011100010011101111101111001111010101111010110";
                    when "01010" => level_vec_out <= "0111111111111111111011100010011101111101111001111010101111010110";
                    when "01011" => level_vec_out <= "0111111111111111111011110010011101111101111001111010101111010110";
                    when "01100" => level_vec_out <= "1111111111111111111011110010011101111101111001111010101111010110";
                    when "01101" => level_vec_out <= "1111111111111111111011110110011101111101111001111010101111010110";
                    when "01110" => level_vec_out <= "1111111111111111111011110110011101111101111001111010101111010110";
                    when "01111" => level_vec_out <= "1111111111111111111011110111011101111101111001111010101111010110";
                    when "10000" => level_vec_out <= "1111111111111111111011110111011101111101111001111110101111010110";
                    when "10001" => level_vec_out <= "1111111111111111111011110111011101111101111001111110101111010110";
                    when "10010" => level_vec_out <= "1111111111111111111011110111011101111101111001111110101111010110";
                    when "10011" => level_vec_out <= "1111111111111111111011110111011101111101111001111110101111010110";
                    when "10100" => level_vec_out <= "1111111111111111111011110111011101111111111001111110101111010110";
                    when "10101" => level_vec_out <= "1111111111111111111011110111111101111111111001111110101111010110";
                    when "10110" => level_vec_out <= "1111111111111111111011110111111101111111111001111110101111010110";
                    when "10111" => level_vec_out <= "1111111111111111111011110111111111111111111111111110101111110110";
                    when "11000" => level_vec_out <= "1111111111111111111011110111111111111111111111111110101111110110";
                    when "11001" => level_vec_out <= "1111111111111111111011110111111111111111111111111110111111110110";
                    when "11010" => level_vec_out <= "1111111111111111111011110111111111111111111111111110111111111110";
                    when "11011" => level_vec_out <= "1111111111111111111011110111111111111111111111111110111111111110";
                    when "11100" => level_vec_out <= "1111111111111111111011111111111111111111111111111110111111111111";
                    when "11101" => level_vec_out <= "1111111111111111111011111111111111111111111111111111111111111111";
                    when "11110" => level_vec_out <= "1111111111111111111011111111111111111111111111111111111111111111";
                    when "11111" => level_vec_out <= "1111111111111111111011111111111111111111111111111111111111111111";
                when others => null;
                end case;
            when others => null;
        end case;
    end process;
end Behavioral;