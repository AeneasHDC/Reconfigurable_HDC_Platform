/**
 * @file level_hvec_gen_hdl.hpp
 * @brief This script generates HDL code for generating high-dimensional LEVEL vectors.
 * It is a novel method; for more information, please refer to our paper.
 *
 * @author Saeid Jamili and Marco Angioli
 * @note Author names are listed in alphabetical order.
 * @email <saeid.jamili@uniroma1.it>
 * @email <marco.angioli@uniroma1.it>
 *
 * @contributors
 *
 * @date Created: 24th July 2023
 * @date Last Updated: 23th August 2023
 *
 * @version 1.0.0
 *
 * @institute Sapienza University of Rome
 * @cite https://doi.org/10.xxxx/yyyyy
 *
 * @section DEPENDENCIES
 * - Dependency1: Description or version details.
 * - Dependency2: Description or version details.
 *
 * @section LICENSE
 * This file is part of the Aeneas HyperCompute Platform.
 *
 * Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 *
 * @section CHANGELOG
 * @version 1.0.0-dev - 23th August 2023
 * - Initial release
 *
 * @todo
 * - Complete level vector generator function
 * - Add training
 *
 * @see
 * -
 * -
 * -
 *
 */

module level_hvec_gen #(parameter int DI_PARALLEL_W_BITS = 64) (
  input logic [2:0] frame_index,
  input logic [4:0] frame_id,
  output logic [DI_PARALLEL_W_BITS-1:0] level_vec_out
);
  always_comb begin
    case (frame_index)
      0:
        case (frame_id)
          0:
            level_vec_out = 64'b1000011101100110111100111000100101000001100010111000000101111110;
          1:
            level_vec_out = 64'b1000011101100110111100111000100101010001100010111100000101111110;
          2:
            level_vec_out = 64'b1000011101100110111100111000100101110001100010111100000101111110;
          3:
            level_vec_out = 64'b1000011101100110111100111000100101110001100010111100000101111110;
          4:
            level_vec_out = 64'b1010011101100110111100111000100101110001100010111100001101111110;
          5:
            level_vec_out = 64'b1010011101100110111100111000100101110011100010111100001101111110;
          6:
            level_vec_out = 64'b1010011101100110111100111000100101110011100010111100001101111110;
          7:
            level_vec_out = 64'b1010011101100110111100111000100101110011100010111100001101111110;
          8:
            level_vec_out = 64'b1110011101100110111100111000100101110011100010111100001101111110;
          9:
            level_vec_out = 64'b1110011101100110111100111000110101110011100011111100001101111110;
          10:
            level_vec_out = 64'b1110011101100110111100111000110111110011100011111100001101111110;
          11:
            level_vec_out = 64'b1110011101100110111101111000110111110011100011111100001101111110;
          12:
            level_vec_out = 64'b1110011101100110111101111000111111110011100011111100001101111110;
          13:
            level_vec_out = 64'b1110011101100110111101111000111111110011100011111101001101111110;
          14:
            level_vec_out = 64'b1110011101100110111101111000111111110011100011111101001101111110;
          15:
            level_vec_out = 64'b1110011101100110111101111000111111110011100011111101101101111110;
          16:
            level_vec_out = 64'b1110011101100110111101111001111111110011100011111101101101111110;
          17:
            level_vec_out = 64'b1110011101100110111101111101111111110011100111111101101101111110;
          18:
            level_vec_out = 64'b1110011111100110111101111101111111110011100111111101101111111110;
          19:
            level_vec_out = 64'b1110111111100110111101111111111111110011100111111101101111111110;
          20:
            level_vec_out = 64'b1110111111100110111101111111111111110011100111111101101111111110;
          21:
            level_vec_out = 64'b1110111111100110111101111111111111110011100111111101101111111110;
          22:
            level_vec_out = 64'b1110111111100110111111111111111111110011100111111101111111111110;
          23:
            level_vec_out = 64'b1110111111100110111111111111111111110011100111111101111111111110;
          24:
            level_vec_out = 64'b1110111111100110111111111111111111110011100111111101111111111110;
          25:
            level_vec_out = 64'b1110111111100111111111111111111111110011100111111101111111111110;
          26:
            level_vec_out = 64'b1110111111110111111111111111111111110011101111111101111111111110;
          27:
            level_vec_out = 64'b1111111111110111111111111111111111110011101111111111111111111110;
          28:
            level_vec_out = 64'b1111111111111111111111111111111111110011101111111111111111111110;
          29:
            level_vec_out = 64'b1111111111111111111111111111111111111011111111111111111111111110;
          30:
            level_vec_out = 64'b1111111111111111111111111111111111111011111111111111111111111110;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        endcase
      1:
        case (frame_id)
          0:
            level_vec_out = 64'b1000111110011111011011001011000011111101111011101110101010110111;
          1:
            level_vec_out = 64'b1000111110011111011011001011001011111101111011101110101010110111;
          2:
            level_vec_out = 64'b1000111110011111011011001011001011111101111011111110101010110111;
          3:
            level_vec_out = 64'b1000111110011111011011101011011111111101111011111110101010110111;
          4:
            level_vec_out = 64'b1000111110011111011011101011011111111101111011111110101010110111;
          5:
            level_vec_out = 64'b1000111110011111011011101011011111111101111011111111101010110111;
          6:
            level_vec_out = 64'b1010111110011111011011101011011111111101111011111111101010110111;
          7:
            level_vec_out = 64'b1011111110011111011011111011011111111101111011111111101010110111;
          8:
            level_vec_out = 64'b1011111110011111011011111011011111111101111011111111101010110111;
          9:
            level_vec_out = 64'b1011111110011111011011111011011111111101111011111111101010110111;
          10:
            level_vec_out = 64'b1011111110011111011011111011011111111101111011111111101010110111;
          11:
            level_vec_out = 64'b1011111110111111011011111011011111111101111011111111101010110111;
          12:
            level_vec_out = 64'b1011111111111111011011111011011111111101111011111111101010110111;
          13:
            level_vec_out = 64'b1111111111111111011011111011011111111101111011111111101010110111;
          14:
            level_vec_out = 64'b1111111111111111011011111011011111111101111011111111101010110111;
          15:
            level_vec_out = 64'b1111111111111111011011111011111111111101111011111111101010110111;
          16:
            level_vec_out = 64'b1111111111111111011011111011111111111101111011111111101010110111;
          17:
            level_vec_out = 64'b1111111111111111011011111011111111111101111011111111101010110111;
          18:
            level_vec_out = 64'b1111111111111111011011111011111111111101111011111111101010110111;
          19:
            level_vec_out = 64'b1111111111111111011011111011111111111101111011111111101010110111;
          20:
            level_vec_out = 64'b1111111111111111011011111011111111111111111011111111101010110111;
          21:
            level_vec_out = 64'b1111111111111111011011111011111111111111111011111111111010110111;
          22:
            level_vec_out = 64'b1111111111111111011011111011111111111111111011111111111011110111;
          23:
            level_vec_out = 64'b1111111111111111011011111011111111111111111011111111111011110111;
          24:
            level_vec_out = 64'b1111111111111111011011111011111111111111111011111111111111110111;
          25:
            level_vec_out = 64'b1111111111111111111111111011111111111111111011111111111111111111;
          26:
            level_vec_out = 64'b1111111111111111111111111011111111111111111011111111111111111111;
          27:
            level_vec_out = 64'b1111111111111111111111111011111111111111111011111111111111111111;
          28:
            level_vec_out = 64'b1111111111111111111111111011111111111111111011111111111111111111;
          29:
            level_vec_out = 64'b1111111111111111111111111011111111111111111011111111111111111111;
          30:
            level_vec_out = 64'b1111111111111111111111111011111111111111111011111111111111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111011111111111111111011111111111111111111;
        endcase
      2:
        case (frame_id)
          0:
            level_vec_out = 64'b1100000000001101011111111101111110001100100010110110011110010101;
          1:
            level_vec_out = 64'b1100000000001111011111111101111110001100100010110110011110010101;
          2:
            level_vec_out = 64'b1100000000001111011111111101111110001100100010110110011110010101;
          3:
            level_vec_out = 64'b1100000000001111011111111101111110001110100010111110011110010101;
          4:
            level_vec_out = 64'b1100000000001111011111111101111110001110100010111110011110010101;
          5:
            level_vec_out = 64'b1100000000001111011111111101111110001110100010111110011110010101;
          6:
            level_vec_out = 64'b1100000000001111011111111101111110001110100010111111111110010101;
          7:
            level_vec_out = 64'b1100000000001111011111111101111110001110100010111111111110010101;
          8:
            level_vec_out = 64'b1100100000001111011111111101111110001110100010111111111110110101;
          9:
            level_vec_out = 64'b1100100000001111011111111101111110001110100010111111111110110101;
          10:
            level_vec_out = 64'b1100100000001111011111111101111110001110100010111111111110110101;
          11:
            level_vec_out = 64'b1100100000001111011111111101111110001110100010111111111110110101;
          12:
            level_vec_out = 64'b1101100000001111011111111101111110001110100010111111111110110101;
          13:
            level_vec_out = 64'b1101101000001111011111111101111110001110110010111111111110110101;
          14:
            level_vec_out = 64'b1101101000001111011111111101111110001110110010111111111110110111;
          15:
            level_vec_out = 64'b1101101000101111011111111101111110001110110010111111111110110111;
          16:
            level_vec_out = 64'b1101101000101111011111111101111110001110110110111111111110110111;
          17:
            level_vec_out = 64'b1101101000101111011111111101111110001110110110111111111110110111;
          18:
            level_vec_out = 64'b1101101000101111011111111101111111001110110110111111111110110111;
          19:
            level_vec_out = 64'b1101101010111111011111111101111111001110110110111111111110110111;
          20:
            level_vec_out = 64'b1101101010111111011111111101111111001110110110111111111110110111;
          21:
            level_vec_out = 64'b1101111010111111011111111101111111001110110110111111111110110111;
          22:
            level_vec_out = 64'b1101111010111111011111111101111111001110110110111111111110111111;
          23:
            level_vec_out = 64'b1101111110111111011111111101111111001110110110111111111110111111;
          24:
            level_vec_out = 64'b1101111110111111011111111101111111001110110110111111111110111111;
          25:
            level_vec_out = 64'b1101111110111111011111111101111111001110110110111111111110111111;
          26:
            level_vec_out = 64'b1101111111111111011111111101111111011110110110111111111110111111;
          27:
            level_vec_out = 64'b1111111111111111011111111101111111011110110110111111111110111111;
          28:
            level_vec_out = 64'b1111111111111111111111111101111111011110110111111111111111111111;
          29:
            level_vec_out = 64'b1111111111111111111111111101111111011111110111111111111111111111;
          30:
            level_vec_out = 64'b1111111111111111111111111111111111011111110111111111111111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111011111110111111111111111111111;
        endcase
      3:
        case (frame_id)
          0:
            level_vec_out = 64'b1000101000001111001000000001101011010100001110010010110000100111;
          1:
            level_vec_out = 64'b1000101000001111001010000001101011110100001110010010110000100111;
          2:
            level_vec_out = 64'b1000101000001111001010000001101011110100001110010010110000100111;
          3:
            level_vec_out = 64'b1000101000001111001010000001101011110100001110010010110000100111;
          4:
            level_vec_out = 64'b1100101010001111001010100001101011110100001110010010110000100111;
          5:
            level_vec_out = 64'b1100101010001111001010100101101011110100001110010010110000100111;
          6:
            level_vec_out = 64'b1100101010001111001010100101101011110100011110010010110000100111;
          7:
            level_vec_out = 64'b1100101010001111101010100101101011110100011110010010111000100111;
          8:
            level_vec_out = 64'b1100101010001111101010100101101011110100011110010010111000100111;
          9:
            level_vec_out = 64'b1100101010001111101010100101101011110100011110010010111000100111;
          10:
            level_vec_out = 64'b1100101010001111101010110101101011110100011110010010111100100111;
          11:
            level_vec_out = 64'b1100101010001111101010110101101111110100011110010010111100100111;
          12:
            level_vec_out = 64'b1100101010001111101010110101101111110100011110010010111100100111;
          13:
            level_vec_out = 64'b1100101010001111101010110101101111110100011110010110111110100111;
          14:
            level_vec_out = 64'b1100101010001111101011110101101111110100011110010110111110100111;
          15:
            level_vec_out = 64'b1100101010001111101011110101101111110100011110010110111111100111;
          16:
            level_vec_out = 64'b1100101010001111101011110101101111110100011110010110111111100111;
          17:
            level_vec_out = 64'b1100101010001111101011111101101111110100011110010110111111100111;
          18:
            level_vec_out = 64'b1100101010001111101011111101101111110110011110010110111111100111;
          19:
            level_vec_out = 64'b1100101010001111101011111101101111110110011110010110111111100111;
          20:
            level_vec_out = 64'b1110101010001111101111111101101111110110011110010110111111110111;
          21:
            level_vec_out = 64'b1110101010001111101111111101101111110110011110110110111111111111;
          22:
            level_vec_out = 64'b1110101010001111101111111101101111110110011110110110111111111111;
          23:
            level_vec_out = 64'b1110101011001111101111111101101111110110011110110110111111111111;
          24:
            level_vec_out = 64'b1110111011001111101111111101101111110110011111110110111111111111;
          25:
            level_vec_out = 64'b1110111011001111101111111111101111110110011111110110111111111111;
          26:
            level_vec_out = 64'b1110111011001111111111111111101111110110011111110110111111111111;
          27:
            level_vec_out = 64'b1110111111101111111111111111101111110110011111110110111111111111;
          28:
            level_vec_out = 64'b1110111111101111111111111111101111110111011111110110111111111111;
          29:
            level_vec_out = 64'b1110111111101111111111111111101111110111011111110110111111111111;
          30:
            level_vec_out = 64'b1111111111101111111111111111101111111111011111110111111111111111;
          31:
            level_vec_out = 64'b1111111111101111111111111111111111111111011111110111111111111111;
        endcase
      4:
        case (frame_id)
          0:
            level_vec_out = 64'b1001010010000001000001110010000010010010100110001010001001001010;
          1:
            level_vec_out = 64'b1001010010010001000001110010000010010010100110001010001001101010;
          2:
            level_vec_out = 64'b1001010010010001100001110010000010010010100110001010001001111010;
          3:
            level_vec_out = 64'b1001010010010001100001110010000010010010100110001010001001111010;
          4:
            level_vec_out = 64'b1001010010010001100001110010000010010010100110001010001001111010;
          5:
            level_vec_out = 64'b1001010010010101100001110010000010010010100111001110001001111010;
          6:
            level_vec_out = 64'b1001010010010101100001110010000010010010100111001110001011111010;
          7:
            level_vec_out = 64'b1001010010010101100001110010000010010010100111001110001011111010;
          8:
            level_vec_out = 64'b1001010010010101100001110010000010110010100111011110001011111010;
          9:
            level_vec_out = 64'b1001010010010101100101110010000010110010100111111110001011111010;
          10:
            level_vec_out = 64'b1001011010010101100101110010000010110010100111111110001111111010;
          11:
            level_vec_out = 64'b1001011010010101100111110010000010110011100111111110001111111010;
          12:
            level_vec_out = 64'b1001011010010111100111110010010010110011100111111110101111111010;
          13:
            level_vec_out = 64'b1001011010010111100111110010010010110011100111111110101111111010;
          14:
            level_vec_out = 64'b1001011010110111100111110011010010110011100111111110101111111010;
          15:
            level_vec_out = 64'b1001011011110111100111111011010010110011100111111110101111111010;
          16:
            level_vec_out = 64'b1001011011110111100111111011010010110011100111111110101111111010;
          17:
            level_vec_out = 64'b1001011011110111100111111011010010110011100111111110101111111010;
          18:
            level_vec_out = 64'b1001011111110111100111111011010010110111100111111110101111111010;
          19:
            level_vec_out = 64'b1001011111110111100111111011011010110111100111111110101111111110;
          20:
            level_vec_out = 64'b1001011111110111100111111011111010110111100111111110101111111110;
          21:
            level_vec_out = 64'b1001011111110111100111111011111010110111100111111110101111111110;
          22:
            level_vec_out = 64'b1001011111110111101111111011111010110111100111111110101111111110;
          23:
            level_vec_out = 64'b1001011111110111101111111111111010110111100111111110101111111110;
          24:
            level_vec_out = 64'b1001011111110111111111111111111010111111100111111110101111111110;
          25:
            level_vec_out = 64'b1001011111110111111111111111111011111111100111111110101111111111;
          26:
            level_vec_out = 64'b1001011111110111111111111111111111111111100111111111101111111111;
          27:
            level_vec_out = 64'b1001011111110111111111111111111111111111101111111111101111111111;
          28:
            level_vec_out = 64'b1001011111110111111111111111111111111111111111111111101111111111;
          29:
            level_vec_out = 64'b1011011111111111111111111111111111111111111111111111111111111111;
          30:
            level_vec_out = 64'b1011111111111111111111111111111111111111111111111111111111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        endcase
      5:
        case (frame_id)
          0:
            level_vec_out = 64'b1110000000101001101100011010101111110001111010001101111000001001;
          1:
            level_vec_out = 64'b1110000000101001101100011010101111110001111010001101111000001001;
          2:
            level_vec_out = 64'b1110000000101001101101011010101111110001111010001101111000001001;
          3:
            level_vec_out = 64'b1110000000101001101101011110101111110001111010001101111000001001;
          4:
            level_vec_out = 64'b1110000000101001111101011110101111110001111010001101111000001001;
          5:
            level_vec_out = 64'b1110000000101001111101011110101111110001111010001101111100001001;
          6:
            level_vec_out = 64'b1110100000101001111101011110101111110001111010001101111100101001;
          7:
            level_vec_out = 64'b1110100010101001111101011110101111110101111010001101111100101001;
          8:
            level_vec_out = 64'b1110101010101001111101011110101111110111111110001101111100101001;
          9:
            level_vec_out = 64'b1110101010101001111101011110101111110111111110011101111100101001;
          10:
            level_vec_out = 64'b1110101010101001111101011110101111110111111110011111111100101001;
          11:
            level_vec_out = 64'b1110101010101101111101011110101111111111111110011111111100101001;
          12:
            level_vec_out = 64'b1110101010101101111101011110101111111111111110011111111100101001;
          13:
            level_vec_out = 64'b1110101010101101111101011110101111111111111110011111111100101001;
          14:
            level_vec_out = 64'b1110101010101101111101111110101111111111111110011111111100101001;
          15:
            level_vec_out = 64'b1110101010101101111101111110101111111111111111011111111100101001;
          16:
            level_vec_out = 64'b1110101011101101111111111110101111111111111111011111111100101001;
          17:
            level_vec_out = 64'b1110101011101101111111111110101111111111111111011111111100101001;
          18:
            level_vec_out = 64'b1110101011101101111111111110101111111111111111111111111100101001;
          19:
            level_vec_out = 64'b1110101011101101111111111110101111111111111111111111111101101001;
          20:
            level_vec_out = 64'b1110101011101111111111111110101111111111111111111111111101101001;
          21:
            level_vec_out = 64'b1110101011101111111111111110101111111111111111111111111101101001;
          22:
            level_vec_out = 64'b1110101011101111111111111110111111111111111111111111111101101001;
          23:
            level_vec_out = 64'b1111101111101111111111111110111111111111111111111111111101101001;
          24:
            level_vec_out = 64'b1111101111101111111111111111111111111111111111111111111101101001;
          25:
            level_vec_out = 64'b1111101111101111111111111111111111111111111111111111111101101001;
          26:
            level_vec_out = 64'b1111101111101111111111111111111111111111111111111111111101101101;
          27:
            level_vec_out = 64'b1111101111101111111111111111111111111111111111111111111101101101;
          28:
            level_vec_out = 64'b1111101111111111111111111111111111111111111111111111111111101101;
          29:
            level_vec_out = 64'b1111101111111111111111111111111111111111111111111111111111101101;
          30:
            level_vec_out = 64'b1111101111111111111111111111111111111111111111111111111111111101;
          31:
            level_vec_out = 64'b1111101111111111111111111111111111111111111111111111111111111111;
        endcase
      6:
        case (frame_id)
          0:
            level_vec_out = 64'b0000011101101100111101011001100000010111111100000101111100100110;
          1:
            level_vec_out = 64'b0000011101101100111101011001100000010111111100000101111100100110;
          2:
            level_vec_out = 64'b0001011101101100111101011001100000010111111100000101111100100110;
          3:
            level_vec_out = 64'b0001011101101100111101011001100000110111111100000101111100100110;
          4:
            level_vec_out = 64'b0001011101101100111101011011100000110111111100100101111100100110;
          5:
            level_vec_out = 64'b0001011101101100111101011011100000110111111100100101111100100110;
          6:
            level_vec_out = 64'b0001011101101100111101011011100000110111111100100101111100100110;
          7:
            level_vec_out = 64'b1001011101101100111101011011100000110111111100100101111101100110;
          8:
            level_vec_out = 64'b1001011101101100111101011011100000110111111100100101111101100110;
          9:
            level_vec_out = 64'b1001011101101100111101011011100000110111111100100101111101110110;
          10:
            level_vec_out = 64'b1001011101101101111101011011100000110111111100100101111101110110;
          11:
            level_vec_out = 64'b1001011101101101111101011011110000110111111100100101111101110110;
          12:
            level_vec_out = 64'b1001011101101101111101011011110001110111111100100101111101110110;
          13:
            level_vec_out = 64'b1001011101101101111101011011110001110111111100100101111101111110;
          14:
            level_vec_out = 64'b1001011101101101111101011011110001110111111100110101111101111110;
          15:
            level_vec_out = 64'b1001011101101101111101011011110001110111111101110101111101111110;
          16:
            level_vec_out = 64'b1001011101101111111101011011110001110111111101110101111101111110;
          17:
            level_vec_out = 64'b1001111101101111111101011011110011110111111101110101111101111111;
          18:
            level_vec_out = 64'b1001111101101111111101011011110011110111111101110101111101111111;
          19:
            level_vec_out = 64'b1001111101101111111101011011110011110111111101111101111101111111;
          20:
            level_vec_out = 64'b1001111101101111111101011011110011111111111101111101111101111111;
          21:
            level_vec_out = 64'b1001111101111111111111011011110011111111111111111101111101111111;
          22:
            level_vec_out = 64'b1001111111111111111111011011110011111111111111111101111101111111;
          23:
            level_vec_out = 64'b1011111111111111111111011011110011111111111111111101111101111111;
          24:
            level_vec_out = 64'b1011111111111111111111011011110011111111111111111111111111111111;
          25:
            level_vec_out = 64'b1011111111111111111111011011110011111111111111111111111111111111;
          26:
            level_vec_out = 64'b1011111111111111111111011011110011111111111111111111111111111111;
          27:
            level_vec_out = 64'b1011111111111111111111011111110011111111111111111111111111111111;
          28:
            level_vec_out = 64'b1011111111111111111111011111110011111111111111111111111111111111;
          29:
            level_vec_out = 64'b1011111111111111111111011111111011111111111111111111111111111111;
          30:
            level_vec_out = 64'b1011111111111111111111011111111011111111111111111111111111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        endcase
      7:
        case (frame_id)
          0:
            level_vec_out = 64'b0000101111100111010111010011111000001011011001111110101010001110;
          1:
            level_vec_out = 64'b0000101111100111010111010011111000001011011001111110101010001110;
          2:
            level_vec_out = 64'b0000101111100111010111010011111000001111111001111110101010001110;
          3:
            level_vec_out = 64'b0000101111100111010111010011111000001111111001111110101010101110;
          4:
            level_vec_out = 64'b0000101111100111010111010011111000001111111001111110101010101110;
          5:
            level_vec_out = 64'b0000101111100111010111010011111000001111111101111110101010101110;
          6:
            level_vec_out = 64'b0000101111100111010111010011111000001111111101111110101011101110;
          7:
            level_vec_out = 64'b0000101111100111010111010011111000001111111101111110101011101110;
          8:
            level_vec_out = 64'b0000101111100111010111010011111000001111111101111110101011101110;
          9:
            level_vec_out = 64'b0000101111100111010111010011111000001111111101111110101111101111;
          10:
            level_vec_out = 64'b0000101111100111010111010011111000001111111101111110111111101111;
          11:
            level_vec_out = 64'b0000101111100111010111010011111000001111111101111110111111101111;
          12:
            level_vec_out = 64'b0001101111100111010111010011111000001111111101111110111111101111;
          13:
            level_vec_out = 64'b1001101111100111010111010011111000001111111101111110111111101111;
          14:
            level_vec_out = 64'b1001101111100111010111011111111000001111111101111110111111101111;
          15:
            level_vec_out = 64'b1001101111100111010111011111111000001111111101111110111111101111;
          16:
            level_vec_out = 64'b1001101111100111010111011111111011001111111101111111111111101111;
          17:
            level_vec_out = 64'b1001101111111111010111011111111011001111111101111111111111101111;
          18:
            level_vec_out = 64'b1001101111111111010111011111111011001111111111111111111111101111;
          19:
            level_vec_out = 64'b1001101111111111010111011111111011001111111111111111111111101111;
          20:
            level_vec_out = 64'b1101101111111111010111011111111011001111111111111111111111101111;
          21:
            level_vec_out = 64'b1101101111111111010111011111111111001111111111111111111111101111;
          22:
            level_vec_out = 64'b1101111111111111010111011111111111001111111111111111111111101111;
          23:
            level_vec_out = 64'b1111111111111111110111011111111111001111111111111111111111101111;
          24:
            level_vec_out = 64'b1111111111111111110111011111111111001111111111111111111111101111;
          25:
            level_vec_out = 64'b1111111111111111110111011111111111101111111111111111111111101111;
          26:
            level_vec_out = 64'b1111111111111111110111011111111111101111111111111111111111101111;
          27:
            level_vec_out = 64'b1111111111111111111111011111111111101111111111111111111111101111;
          28:
            level_vec_out = 64'b1111111111111111111111011111111111101111111111111111111111101111;
          29:
            level_vec_out = 64'b1111111111111111111111111111111111101111111111111111111111101111;
          30:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
          31:
            level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        endcase
    endcase
  end
endmodule