/**
 * @file level_hvec_gen_hdl.hpp
 * @brief This script generates HDL code for generating high-dimensional LEVEL vectors.
 * It is a novel method; for more information, please refer to our paper.
 *
 * @author Saeid Jamili and Marco Angioli
 * @note Author names are listed in alphabetical order.
 * @email <saeid.jamili@uniroma1.it>
 * @email <marco.angioli@uniroma1.it>
 *
 * @contributors
 *
 * @date Created: 24th July 2023
 * @date Last Updated: 23th August 2023
 *
 * @version 1.0.0
 *
 * @institute Sapienza University of Rome
 * @cite https://doi.org/10.xxxx/yyyyy
 *
 * @section DEPENDENCIES
 * - Dependency1: Description or version details.
 * - Dependency2: Description or version details.
 *
 * @section LICENSE
 * This file is part of the Aeneas HyperCompute Platform.
 *
 * Licensed under the MIT License. See the LICENSE file in the project root for full license details.
 *
 * @section CHANGELOG
 * @version 1.0.0-dev - 23th August 2023
 * - Initial release
 *
 * @todo
 * - Complete level vector generator function
 * - Add training
 *
 * @see
 * -
 * -
 * -
 *
 */

module level_vec_gen (
    output reg [63:0] level_vec_out,
    input [2:0] frame_index,
    input [4:0] frame_id
);
    always @(*) begin
        // Update this function to match your requirements
        case (frame_index)
            0: begin
                case (frame_id)
                    0: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    1: level_vec_out = 64'b1111111111111111000000000000000000000000000000000000000000000000;
                    2: level_vec_out = 64'b1111111111111111111111110000000000000000000000000000000000000000;
                    3: level_vec_out = 64'b1111111111111111111111111111111100000000000000000000000000000000;
                    4: level_vec_out = 64'b1111111111111111111111111111111111111111000000000000000000000000;
                    5: level_vec_out = 64'b1111111111111111111111111111111111111111111111110000000000000000;
                    6: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111100000000;
                    7: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    8: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    9: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    10: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    11: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    12: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    13: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    14: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    15: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    16: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    17: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    18: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    19: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    20: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    21: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    22: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    23: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    24: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    25: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    26: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    27: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    28: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    29: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    30: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    31: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                endcase
            end
            1: begin
                case (frame_id)
                    0: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    1: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    2: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    3: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    4: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    5: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    6: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    7: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    8: level_vec_out = 64'b1111111100000000000000000000000000000000000000000000000000000000;
                    9: level_vec_out = 64'b1111111111111111000000000000000000000000000000000000000000000000;
                    10: level_vec_out = 64'b1111111111111111111111110000000000000000000000000000000000000000;
                    11: level_vec_out = 64'b1111111111111111111111111111111100000000000000000000000000000000;
                    12: level_vec_out = 64'b1111111111111111111111111111111111111111000000000000000000000000;
                    13: level_vec_out = 64'b1111111111111111111111111111111111111111111111110000000000000000;
                    14: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111100000000;
                    15: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    16: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    17: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    18: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    19: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    20: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    21: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    22: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    23: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    24: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    25: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    26: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    27: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    28: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    29: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    30: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    31: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                endcase
            end
            2: begin
                case (frame_id)
                    0: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    1: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    2: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    3: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    4: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    5: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    6: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    7: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    8: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    9: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    10: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    11: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    12: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    13: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    14: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    15: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    16: level_vec_out = 64'b1111111100000000000000000000000000000000000000000000000000000000;
                    17: level_vec_out = 64'b1111111111111111000000000000000000000000000000000000000000000000;
                    18: level_vec_out = 64'b1111111111111111111111110000000000000000000000000000000000000000;
                    19: level_vec_out = 64'b1111111111111111111111111111111100000000000000000000000000000000;
                    20: level_vec_out = 64'b1111111111111111111111111111111111111111000000000000000000000000;
                    21: level_vec_out = 64'b1111111111111111111111111111111111111111111111110000000000000000;
                    22: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111100000000;
                    23: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    24: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    25: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    26: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    27: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    28: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    29: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    30: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                    31: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                endcase
            end
            3: begin
                case (frame_id)
                    0: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    1: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    2: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    3: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    4: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    5: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    6: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    7: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    8: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    9: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    10: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    11: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    12: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    13: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    14: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    15: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    16: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    17: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    18: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    19: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    20: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    21: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    22: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    23: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    24: level_vec_out = 64'b1111111100000000000000000000000000000000000000000000000000000000;
                    25: level_vec_out = 64'b1111111111111111000000000000000000000000000000000000000000000000;
                    26: level_vec_out = 64'b1111111111111111111111110000000000000000000000000000000000000000;
                    27: level_vec_out = 64'b1111111111111111111111111111111100000000000000000000000000000000;
                    28: level_vec_out = 64'b1111111111111111111111111111111111111111000000000000000000000000;
                    29: level_vec_out = 64'b1111111111111111111111111111111111111111111111110000000000000000;
                    30: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111100000000;
                    31: level_vec_out = 64'b1111111111111111111111111111111111111111111111111111111111111111;
                endcase
            end
            4: begin
                case (frame_id)
                    0: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    1: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    2: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    3: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    4: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    5: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    6: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    7: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    8: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    9: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    10: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    11: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    12: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    13: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    14: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    15: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    16: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    17: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    18: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    19: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    20: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    21: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    22: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    23: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    24: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    25: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    26: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    27: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    28: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    29: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    30: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    31: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                endcase
            end
            5: begin
                case (frame_id)
                    0: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    1: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    2: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    3: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    4: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    5: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    6: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    7: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    8: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    9: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    10: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    11: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    12: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    13: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    14: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    15: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    16: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    17: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    18: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    19: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    20: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    21: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    22: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    23: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    24: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    25: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    26: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    27: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    28: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    29: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    30: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    31: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                endcase
            end
            6: begin
                case (frame_id)
                    0: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    1: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    2: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    3: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    4: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    5: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    6: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    7: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    8: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    9: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    10: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    11: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    12: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    13: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    14: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    15: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    16: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    17: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    18: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    19: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    20: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    21: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    22: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    23: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    24: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    25: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    26: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    27: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    28: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    29: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    30: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    31: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                endcase
            end
            7: begin
                case (frame_id)
                    0: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    1: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    2: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    3: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    4: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    5: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    6: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    7: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    8: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    9: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    10: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    11: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    12: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    13: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    14: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    15: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    16: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    17: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    18: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    19: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    20: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    21: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    22: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    23: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    24: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    25: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    26: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    27: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    28: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    29: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    30: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                    31: level_vec_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;
                endcase
            end
        endcase
    end
endmodule